library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity RAM_VIDEO is
  port ( 
    clk  : in    std_logic;   
    addr : in    unsigned (16 downto 0); 
    do   : out   unsigned(23 downto 0)
    );
end RAM_VIDEO;

architecture Behavioral of RAM_VIDEO is
  subtype mot is unsigned( 23 downto 0 );
  type zone_memoire is array (natural range 0 to 640*480/4-1) of mot;
  signal ROM: zone_memoire :=(
   0 => x"ffffff",
   1 => x"ffffff",
   2 => x"ffffff",
   3 => x"ffffff",
   4 => x"ffffff",
   5 => x"ffffff",
   6 => x"ffffff",
   7 => x"ffffff",
   8 => x"ffffff",
   9 => x"ffffff",
   10 => x"ffffff",
   11 => x"ffffff",
   12 => x"ffffff",
   13 => x"ffffff",
   14 => x"ffffff",
   15 => x"ffffff",
   16 => x"ffffff",
   17 => x"ffffff",
   18 => x"ffffff",
   19 => x"ffffff",
   20 => x"ffffff",
   21 => x"ffffff",
   22 => x"ffffff",
   23 => x"ffffff",
   24 => x"ffffff",
   25 => x"ffffff",
   26 => x"ffffff",
   27 => x"ffffff",
   28 => x"ffffff",
   29 => x"ffffff",
   30 => x"ffffff",
   31 => x"ffffff",
   32 => x"ffffff",
   33 => x"ffffff",
   34 => x"ffffff",
   35 => x"ffffff",
   36 => x"ffffff",
   37 => x"ffffff",
   38 => x"ffffff",
   39 => x"ffffff",
   40 => x"ffffff",
   41 => x"ffffff",
   42 => x"ffffff",
   43 => x"ffffff",
   44 => x"ffffff",
   45 => x"ffffff",
   46 => x"ffffff",
   47 => x"ffffff",
   48 => x"ffffff",
   49 => x"ffffff",
   50 => x"ffffff",
   51 => x"ffffff",
   52 => x"ffffff",
   53 => x"ffffff",
   54 => x"ffffff",
   55 => x"ffffff",
   56 => x"ffffff",
   57 => x"ffffff",
   58 => x"ffffff",
   59 => x"ffffff",
   60 => x"ffffff",
   61 => x"ffffff",
   62 => x"ffffff",
   63 => x"ffffff",
   64 => x"ffffff",
   65 => x"ffffff",
   66 => x"ffffff",
   67 => x"ffffff",
   68 => x"ffffff",
   69 => x"ffffff",
   70 => x"ffffff",
   71 => x"ffffff",
   72 => x"ffffff",
   73 => x"ffffff",
   74 => x"ffffff",
   75 => x"ffffff",
   76 => x"ffffff",
   77 => x"ffffff",
   78 => x"ffffff",
   79 => x"ffffff",
   80 => x"ffffff",
   81 => x"ffffff",
   82 => x"ffffff",
   83 => x"ffffff",
   84 => x"ffffff",
   85 => x"ffffff",
   86 => x"ffffff",
   87 => x"ffffff",
   88 => x"ffffff",
   89 => x"ffffff",
   90 => x"ffffff",
   91 => x"ffffff",
   92 => x"ffffff",
   93 => x"ffffff",
   94 => x"ffffff",
   95 => x"ffffff",
   96 => x"ffffff",
   97 => x"ffffff",
   98 => x"ffffff",
   99 => x"ffffff",
   100 => x"ffffff",
   101 => x"ffffff",
   102 => x"ffffff",
   103 => x"ffffff",
   104 => x"ffffff",
   105 => x"ffffff",
   106 => x"ffffff",
   107 => x"ffffff",
   108 => x"ffffff",
   109 => x"ffffff",
   110 => x"ffffff",
   111 => x"fffaaa",
   112 => x"aaaaaa",
   113 => x"aaaaaa",
   114 => x"aaaaaa",
   115 => x"aaaaaa",
   116 => x"aaaaaa",
   117 => x"aaaaaa",
   118 => x"aaaaaa",
   119 => x"aaaaaa",
   120 => x"aaaaaa",
   121 => x"aaaaaa",
   122 => x"aaaaaa",
   123 => x"aaaaaa",
   124 => x"aaaaaa",
   125 => x"a95555",
   126 => x"555555",
   127 => x"555555",
   128 => x"555555",
   129 => x"555555",
   130 => x"555555",
   131 => x"555555",
   132 => x"555555",
   133 => x"555555",
   134 => x"555555",
   135 => x"555555",
   136 => x"555555",
   137 => x"555555",
   138 => x"555555",
   139 => x"555555",
   140 => x"555555",
   141 => x"555555",
   142 => x"555555",
   143 => x"555555",
   144 => x"555555",
   145 => x"555555",
   146 => x"555555",
   147 => x"555555",
   148 => x"540000",
   149 => x"000000",
   150 => x"000000",
   151 => x"000000",
   152 => x"000000",
   153 => x"000000",
   154 => x"000000",
   155 => x"000000",
   156 => x"02afff",
   157 => x"ffffff",
   158 => x"ffffff",
   159 => x"ffffff",
   160 => x"ffffff",
   161 => x"ffffff",
   162 => x"ffffff",
   163 => x"ffffff",
   164 => x"ffffff",
   165 => x"ffffff",
   166 => x"ffffff",
   167 => x"ffffff",
   168 => x"ffffff",
   169 => x"ffffff",
   170 => x"ffffff",
   171 => x"ffffff",
   172 => x"ffffff",
   173 => x"ffffff",
   174 => x"ffffff",
   175 => x"ffffff",
   176 => x"ffffff",
   177 => x"ffffff",
   178 => x"ffffff",
   179 => x"ffffff",
   180 => x"ffffff",
   181 => x"ffffff",
   182 => x"ffffff",
   183 => x"ffffff",
   184 => x"ffffff",
   185 => x"ffffff",
   186 => x"ffffff",
   187 => x"ffffff",
   188 => x"ffffff",
   189 => x"ffffff",
   190 => x"ffffff",
   191 => x"ffffff",
   192 => x"ffffff",
   193 => x"ffffff",
   194 => x"ffffff",
   195 => x"ffffff",
   196 => x"ffffff",
   197 => x"ffffff",
   198 => x"ffffff",
   199 => x"ffffff",
   200 => x"ffffff",
   201 => x"ffffff",
   202 => x"ffffff",
   203 => x"ffffff",
   204 => x"ffffff",
   205 => x"ffffff",
   206 => x"ffffff",
   207 => x"ffffff",
   208 => x"ffffff",
   209 => x"ffffff",
   210 => x"ffffff",
   211 => x"ffffff",
   212 => x"ffffff",
   213 => x"ffffff",
   214 => x"ffffff",
   215 => x"ffffff",
   216 => x"ffffff",
   217 => x"ffffff",
   218 => x"ffffff",
   219 => x"ffffff",
   220 => x"ffffff",
   221 => x"ffffff",
   222 => x"ffffff",
   223 => x"ffffff",
   224 => x"ffffff",
   225 => x"ffffff",
   226 => x"ffffff",
   227 => x"ffffff",
   228 => x"ffffff",
   229 => x"ffffff",
   230 => x"ffffff",
   231 => x"ffffff",
   232 => x"ffffff",
   233 => x"ffffff",
   234 => x"ffffff",
   235 => x"ffffff",
   236 => x"ffffff",
   237 => x"ffffff",
   238 => x"ffffff",
   239 => x"ffffff",
   240 => x"ffffff",
   241 => x"ffffff",
   242 => x"ffffff",
   243 => x"ffffff",
   244 => x"ffffff",
   245 => x"ffffff",
   246 => x"ffffff",
   247 => x"ffffff",
   248 => x"ffffff",
   249 => x"ffffff",
   250 => x"ffffff",
   251 => x"ffffff",
   252 => x"ffffff",
   253 => x"ffffff",
   254 => x"ffffff",
   255 => x"ffffff",
   256 => x"ffffff",
   257 => x"ffffff",
   258 => x"ffffff",
   259 => x"ffffff",
   260 => x"ffffff",
   261 => x"ffffff",
   262 => x"ffffff",
   263 => x"ffffff",
   264 => x"ffffff",
   265 => x"ffffff",
   266 => x"ffffff",
   267 => x"ffffff",
   268 => x"ffffff",
   269 => x"ffffff",
   270 => x"ffffff",
   271 => x"fea555",
   272 => x"555555",
   273 => x"555555",
   274 => x"555555",
   275 => x"555555",
   276 => x"555555",
   277 => x"555555",
   278 => x"555555",
   279 => x"555555",
   280 => x"555555",
   281 => x"555555",
   282 => x"555555",
   283 => x"555555",
   284 => x"56aaaa",
   285 => x"aaaaaa",
   286 => x"aaaaaa",
   287 => x"aaaaaa",
   288 => x"aaaaaa",
   289 => x"aaaaaa",
   290 => x"aaaaaa",
   291 => x"aaaaaa",
   292 => x"aaaaaa",
   293 => x"aaaaaa",
   294 => x"aaaaaa",
   295 => x"aaaaaa",
   296 => x"aaaaaa",
   297 => x"aaaaaa",
   298 => x"aaaaaa",
   299 => x"aaaaaa",
   300 => x"aaaaaa",
   301 => x"aaaaaa",
   302 => x"aaaaaa",
   303 => x"aaaaaa",
   304 => x"aaaaaa",
   305 => x"aaaaaa",
   306 => x"aaaaaa",
   307 => x"aaaaaa",
   308 => x"aaaaaa",
   309 => x"aaaaaa",
   310 => x"abffff",
   311 => x"ffffff",
   312 => x"ffffff",
   313 => x"ffffff",
   314 => x"ffffff",
   315 => x"ffffff",
   316 => x"ffffff",
   317 => x"ffffff",
   318 => x"ffffff",
   319 => x"ffffff",
   320 => x"ffffff",
   321 => x"ffffff",
   322 => x"ffffff",
   323 => x"ffffff",
   324 => x"ffffff",
   325 => x"ffffff",
   326 => x"ffffff",
   327 => x"ffffff",
   328 => x"ffffff",
   329 => x"ffffff",
   330 => x"ffffff",
   331 => x"ffffff",
   332 => x"ffffff",
   333 => x"ffffff",
   334 => x"ffffff",
   335 => x"ffffff",
   336 => x"ffffff",
   337 => x"ffffff",
   338 => x"ffffff",
   339 => x"ffffff",
   340 => x"ffffff",
   341 => x"ffffff",
   342 => x"ffffff",
   343 => x"ffffff",
   344 => x"ffffff",
   345 => x"ffffff",
   346 => x"ffffff",
   347 => x"ffffff",
   348 => x"ffffff",
   349 => x"ffffff",
   350 => x"ffffff",
   351 => x"ffffff",
   352 => x"ffffff",
   353 => x"ffffff",
   354 => x"ffffff",
   355 => x"ffffff",
   356 => x"ffffff",
   357 => x"ffffff",
   358 => x"ffffff",
   359 => x"ffffff",
   360 => x"ffffff",
   361 => x"ffffff",
   362 => x"ffffff",
   363 => x"ffffff",
   364 => x"ffffff",
   365 => x"ffffff",
   366 => x"ffffff",
   367 => x"ffffff",
   368 => x"ffffff",
   369 => x"ffffff",
   370 => x"ffffff",
   371 => x"ffffff",
   372 => x"ffffff",
   373 => x"ffffff",
   374 => x"ffffff",
   375 => x"ffffff",
   376 => x"ffffff",
   377 => x"ffffff",
   378 => x"ffffff",
   379 => x"ffffff",
   380 => x"ffffff",
   381 => x"ffffff",
   382 => x"ffffff",
   383 => x"ffffff",
   384 => x"ffffff",
   385 => x"ffffff",
   386 => x"ffffff",
   387 => x"ffffff",
   388 => x"ffffff",
   389 => x"ffffff",
   390 => x"ffffff",
   391 => x"ffffff",
   392 => x"ffffff",
   393 => x"ffffff",
   394 => x"ffffff",
   395 => x"ffffff",
   396 => x"ffffff",
   397 => x"ffffff",
   398 => x"ffffff",
   399 => x"ffffff",
   400 => x"ffffff",
   401 => x"ffffff",
   402 => x"ffffff",
   403 => x"ffffff",
   404 => x"ffffff",
   405 => x"ffffff",
   406 => x"ffffff",
   407 => x"ffffff",
   408 => x"ffffff",
   409 => x"ffffff",
   410 => x"ffffff",
   411 => x"ffffff",
   412 => x"ffffff",
   413 => x"ffffff",
   414 => x"ffffff",
   415 => x"ffffff",
   416 => x"ffffff",
   417 => x"ffffff",
   418 => x"ffffff",
   419 => x"ffffff",
   420 => x"ffffff",
   421 => x"ffffff",
   422 => x"ffffff",
   423 => x"ffffff",
   424 => x"ffffff",
   425 => x"ffffff",
   426 => x"ffffff",
   427 => x"ffffff",
   428 => x"ffffff",
   429 => x"ffffff",
   430 => x"ffffff",
   431 => x"a95abf",
   432 => x"ffffff",
   433 => x"ffffff",
   434 => x"ffffff",
   435 => x"ffffff",
   436 => x"ffffff",
   437 => x"ffffff",
   438 => x"ffffff",
   439 => x"ffffff",
   440 => x"ffffff",
   441 => x"ffffff",
   442 => x"ffffff",
   443 => x"ffffff",
   444 => x"ffffff",
   445 => x"ffffff",
   446 => x"ffffff",
   447 => x"ffffff",
   448 => x"ffffff",
   449 => x"ffffff",
   450 => x"ffffff",
   451 => x"ffffff",
   452 => x"ffffff",
   453 => x"ffffff",
   454 => x"ffffff",
   455 => x"ffffff",
   456 => x"ffffff",
   457 => x"ffffff",
   458 => x"ffffff",
   459 => x"ffffff",
   460 => x"ffffff",
   461 => x"ffffff",
   462 => x"ffffff",
   463 => x"ffffff",
   464 => x"ffffff",
   465 => x"ffffff",
   466 => x"ffffff",
   467 => x"ffffff",
   468 => x"ffffff",
   469 => x"ffffff",
   470 => x"ffffff",
   471 => x"ffffff",
   472 => x"ffffff",
   473 => x"ffffff",
   474 => x"ffffff",
   475 => x"ffffff",
   476 => x"ffffff",
   477 => x"ffffff",
   478 => x"ffffff",
   479 => x"ffffff",
   480 => x"ffffff",
   481 => x"ffffff",
   482 => x"ffffff",
   483 => x"ffffff",
   484 => x"ffffff",
   485 => x"ffffff",
   486 => x"ffffff",
   487 => x"ffffff",
   488 => x"ffffff",
   489 => x"ffffff",
   490 => x"ffffff",
   491 => x"ffffff",
   492 => x"ffffff",
   493 => x"ffffff",
   494 => x"ffffff",
   495 => x"ffffff",
   496 => x"ffffff",
   497 => x"ffffff",
   498 => x"ffffff",
   499 => x"ffffff",
   500 => x"ffffff",
   501 => x"ffffff",
   502 => x"ffffff",
   503 => x"ffffff",
   504 => x"ffffff",
   505 => x"ffffff",
   506 => x"ffffff",
   507 => x"ffffff",
   508 => x"ffffff",
   509 => x"ffffff",
   510 => x"ffffff",
   511 => x"ffffff",
   512 => x"ffffff",
   513 => x"ffffff",
   514 => x"ffffff",
   515 => x"ffffff",
   516 => x"ffffff",
   517 => x"ffffff",
   518 => x"ffffff",
   519 => x"ffffff",
   520 => x"ffffff",
   521 => x"ffffff",
   522 => x"ffffff",
   523 => x"ffffff",
   524 => x"ffffff",
   525 => x"ffffff",
   526 => x"ffffff",
   527 => x"ffffff",
   528 => x"ffffff",
   529 => x"ffffff",
   530 => x"ffffff",
   531 => x"ffffff",
   532 => x"ffffff",
   533 => x"ffffff",
   534 => x"ffffff",
   535 => x"ffffff",
   536 => x"ffffff",
   537 => x"ffffff",
   538 => x"ffffff",
   539 => x"ffffff",
   540 => x"ffffff",
   541 => x"ffffff",
   542 => x"ffffff",
   543 => x"ffffff",
   544 => x"ffffff",
   545 => x"ffffff",
   546 => x"ffffff",
   547 => x"ffffff",
   548 => x"ffffff",
   549 => x"ffffff",
   550 => x"ffffff",
   551 => x"ffffff",
   552 => x"ffffff",
   553 => x"ffffff",
   554 => x"ffffff",
   555 => x"ffffff",
   556 => x"ffffff",
   557 => x"ffffff",
   558 => x"ffffff",
   559 => x"ffffff",
   560 => x"ffffff",
   561 => x"ffffff",
   562 => x"ffffff",
   563 => x"ffffff",
   564 => x"ffffff",
   565 => x"ffffff",
   566 => x"ffffff",
   567 => x"ffffff",
   568 => x"ffffff",
   569 => x"ffffff",
   570 => x"ffffff",
   571 => x"ffffff",
   572 => x"ffffff",
   573 => x"ffffff",
   574 => x"ffffff",
   575 => x"ffffff",
   576 => x"ffffff",
   577 => x"ffffff",
   578 => x"ffffff",
   579 => x"ffffff",
   580 => x"ffffff",
   581 => x"ffffff",
   582 => x"ffffff",
   583 => x"ffffff",
   584 => x"ffffff",
   585 => x"ffffff",
   586 => x"ffffff",
   587 => x"ffffff",
   588 => x"ffffff",
   589 => x"ffffff",
   590 => x"ffffea",
   591 => x"56afff",
   592 => x"ffffff",
   593 => x"ffffff",
   594 => x"ffffff",
   595 => x"ffffff",
   596 => x"ffffff",
   597 => x"ffffff",
   598 => x"ffffff",
   599 => x"ffffff",
   600 => x"ffffff",
   601 => x"ffffff",
   602 => x"ffffff",
   603 => x"ffffff",
   604 => x"ffffff",
   605 => x"ffffff",
   606 => x"ffffff",
   607 => x"ffffff",
   608 => x"ffffff",
   609 => x"ffffff",
   610 => x"ffffff",
   611 => x"ffffff",
   612 => x"ffffff",
   613 => x"ffffff",
   614 => x"ffffff",
   615 => x"ffffff",
   616 => x"ffffff",
   617 => x"ffffff",
   618 => x"ffffff",
   619 => x"ffffff",
   620 => x"ffffff",
   621 => x"ffffff",
   622 => x"ffffff",
   623 => x"ffffff",
   624 => x"ffffff",
   625 => x"ffffff",
   626 => x"ffffff",
   627 => x"ffffff",
   628 => x"ffffff",
   629 => x"ffffff",
   630 => x"ffffff",
   631 => x"ffffff",
   632 => x"ffffff",
   633 => x"ffffff",
   634 => x"ffffff",
   635 => x"ffffff",
   636 => x"ffffff",
   637 => x"ffffff",
   638 => x"ffffff",
   639 => x"ffffff",
   640 => x"ffffff",
   641 => x"ffffff",
   642 => x"ffffff",
   643 => x"ffffff",
   644 => x"ffffff",
   645 => x"ffffff",
   646 => x"ffffff",
   647 => x"ffffff",
   648 => x"ffffff",
   649 => x"ffffff",
   650 => x"ffffff",
   651 => x"ffffff",
   652 => x"ffffff",
   653 => x"ffffff",
   654 => x"ffffff",
   655 => x"ffffff",
   656 => x"ffffff",
   657 => x"ffffff",
   658 => x"ffffff",
   659 => x"ffffff",
   660 => x"ffffff",
   661 => x"ffffff",
   662 => x"ffffff",
   663 => x"ffffff",
   664 => x"ffffff",
   665 => x"ffffff",
   666 => x"ffffff",
   667 => x"ffffff",
   668 => x"ffffff",
   669 => x"ffffff",
   670 => x"ffffff",
   671 => x"ffffff",
   672 => x"ffffff",
   673 => x"ffffff",
   674 => x"ffffff",
   675 => x"ffffff",
   676 => x"ffffff",
   677 => x"ffffff",
   678 => x"ffffff",
   679 => x"ffffff",
   680 => x"ffffff",
   681 => x"ffffff",
   682 => x"ffffff",
   683 => x"ffffff",
   684 => x"ffffff",
   685 => x"ffffff",
   686 => x"ffffff",
   687 => x"ffffff",
   688 => x"ffffff",
   689 => x"ffffff",
   690 => x"ffffff",
   691 => x"ffffff",
   692 => x"ffffff",
   693 => x"ffffff",
   694 => x"ffffff",
   695 => x"ffffff",
   696 => x"ffffff",
   697 => x"ffffff",
   698 => x"ffffff",
   699 => x"ffffff",
   700 => x"ffffff",
   701 => x"ffffff",
   702 => x"ffffff",
   703 => x"fffaaa",
   704 => x"555000",
   705 => x"000015",
   706 => x"56aabf",
   707 => x"ffffff",
   708 => x"ffffff",
   709 => x"ffffff",
   710 => x"ffffff",
   711 => x"ffffff",
   712 => x"ffffff",
   713 => x"ffffff",
   714 => x"ffffff",
   715 => x"ffffff",
   716 => x"ffffff",
   717 => x"ffffff",
   718 => x"ffffff",
   719 => x"ffffff",
   720 => x"ffffff",
   721 => x"ffffff",
   722 => x"ffffff",
   723 => x"ffffff",
   724 => x"ffffff",
   725 => x"ffffff",
   726 => x"ffffff",
   727 => x"ffffff",
   728 => x"ffffff",
   729 => x"ffffff",
   730 => x"ffffff",
   731 => x"ffffff",
   732 => x"ffffff",
   733 => x"ffffff",
   734 => x"ffffff",
   735 => x"ffffff",
   736 => x"ffffff",
   737 => x"ffffff",
   738 => x"ffffff",
   739 => x"ffffff",
   740 => x"ffffff",
   741 => x"ffffff",
   742 => x"ffffff",
   743 => x"ffffff",
   744 => x"ffffff",
   745 => x"ffffff",
   746 => x"ffffff",
   747 => x"ffffff",
   748 => x"ffffff",
   749 => x"ffffff",
   750 => x"fffa95",
   751 => x"abffff",
   752 => x"ffffff",
   753 => x"ffffff",
   754 => x"ffffff",
   755 => x"ffffff",
   756 => x"ffffff",
   757 => x"ffffff",
   758 => x"ffffff",
   759 => x"ffffff",
   760 => x"ffffff",
   761 => x"ffffff",
   762 => x"ffffff",
   763 => x"ffffff",
   764 => x"ffffff",
   765 => x"ffffff",
   766 => x"ffffff",
   767 => x"ffffff",
   768 => x"ffffff",
   769 => x"ffffff",
   770 => x"ffffff",
   771 => x"ffffff",
   772 => x"ffffff",
   773 => x"ffffff",
   774 => x"ffffff",
   775 => x"ffffff",
   776 => x"ffffff",
   777 => x"ffffff",
   778 => x"ffffff",
   779 => x"ffffff",
   780 => x"ffffff",
   781 => x"ffffff",
   782 => x"ffffff",
   783 => x"ffffff",
   784 => x"ffffff",
   785 => x"ffffff",
   786 => x"ffffff",
   787 => x"ffffff",
   788 => x"ffffff",
   789 => x"ffffff",
   790 => x"ffffff",
   791 => x"ffffff",
   792 => x"ffffff",
   793 => x"ffffff",
   794 => x"ffffff",
   795 => x"ffffff",
   796 => x"ffffff",
   797 => x"ffffff",
   798 => x"ffffff",
   799 => x"ffffff",
   800 => x"ffffff",
   801 => x"ffffff",
   802 => x"ffffff",
   803 => x"ffffff",
   804 => x"ffffff",
   805 => x"ffffff",
   806 => x"ffffff",
   807 => x"ffffff",
   808 => x"ffffff",
   809 => x"ffffff",
   810 => x"ffffff",
   811 => x"ffffff",
   812 => x"ffffff",
   813 => x"ffffff",
   814 => x"ffffff",
   815 => x"ffffff",
   816 => x"ffffff",
   817 => x"ffffff",
   818 => x"ffffff",
   819 => x"ffffff",
   820 => x"ffffff",
   821 => x"ffffff",
   822 => x"ffffff",
   823 => x"ffffff",
   824 => x"ffffff",
   825 => x"ffffff",
   826 => x"ffffff",
   827 => x"ffffff",
   828 => x"ffffff",
   829 => x"ffffff",
   830 => x"ffffff",
   831 => x"ffffff",
   832 => x"ffffff",
   833 => x"ffffff",
   834 => x"ffffff",
   835 => x"ffffff",
   836 => x"ffffff",
   837 => x"ffffff",
   838 => x"ffffff",
   839 => x"ffffff",
   840 => x"ffffff",
   841 => x"ffffff",
   842 => x"ffffff",
   843 => x"ffffff",
   844 => x"ffffff",
   845 => x"ffffff",
   846 => x"ffffff",
   847 => x"ffffff",
   848 => x"ffffff",
   849 => x"ffffff",
   850 => x"ffffff",
   851 => x"ffffff",
   852 => x"ffffff",
   853 => x"ffffff",
   854 => x"ffffff",
   855 => x"ffffff",
   856 => x"ffffff",
   857 => x"ffffff",
   858 => x"ffffff",
   859 => x"ffffff",
   860 => x"ffffff",
   861 => x"ffffff",
   862 => x"ffffff",
   863 => x"a95000",
   864 => x"000000",
   865 => x"000000",
   866 => x"000015",
   867 => x"57ffff",
   868 => x"ffffff",
   869 => x"ffffff",
   870 => x"ffffff",
   871 => x"ffffff",
   872 => x"ffffff",
   873 => x"ffffff",
   874 => x"ffffff",
   875 => x"ffffff",
   876 => x"ffffff",
   877 => x"ffffff",
   878 => x"ffffff",
   879 => x"ffffff",
   880 => x"ffffff",
   881 => x"ffffff",
   882 => x"ffffff",
   883 => x"ffffff",
   884 => x"ffffff",
   885 => x"ffffff",
   886 => x"ffffff",
   887 => x"ffffff",
   888 => x"ffffff",
   889 => x"ffffff",
   890 => x"ffffff",
   891 => x"ffffff",
   892 => x"ffffff",
   893 => x"ffffff",
   894 => x"ffffff",
   895 => x"ffffff",
   896 => x"ffffff",
   897 => x"ffffff",
   898 => x"ffffff",
   899 => x"ffffff",
   900 => x"ffffff",
   901 => x"ffffff",
   902 => x"ffffff",
   903 => x"ffffff",
   904 => x"ffffff",
   905 => x"ffffff",
   906 => x"ffffff",
   907 => x"ffffff",
   908 => x"ffffff",
   909 => x"ffffff",
   910 => x"fea56a",
   911 => x"ffffff",
   912 => x"ffffff",
   913 => x"ffffff",
   914 => x"ffffff",
   915 => x"ffffff",
   916 => x"ffffff",
   917 => x"ffffff",
   918 => x"ffffff",
   919 => x"ffffff",
   920 => x"ffffff",
   921 => x"ffffff",
   922 => x"ffffff",
   923 => x"ffffff",
   924 => x"ffffff",
   925 => x"ffffff",
   926 => x"ffffff",
   927 => x"ffffff",
   928 => x"ffffff",
   929 => x"ffffff",
   930 => x"ffffff",
   931 => x"ffffff",
   932 => x"ffffff",
   933 => x"ffffff",
   934 => x"ffffff",
   935 => x"ffffff",
   936 => x"ffffff",
   937 => x"ffffff",
   938 => x"ffffff",
   939 => x"ffffff",
   940 => x"ffffff",
   941 => x"ffffff",
   942 => x"ffffff",
   943 => x"ffffff",
   944 => x"ffffff",
   945 => x"ffffff",
   946 => x"ffffff",
   947 => x"ffffff",
   948 => x"ffffff",
   949 => x"ffffff",
   950 => x"ffffff",
   951 => x"ffffff",
   952 => x"ffffff",
   953 => x"ffffff",
   954 => x"ffffff",
   955 => x"ffffff",
   956 => x"ffffff",
   957 => x"ffffff",
   958 => x"ffffff",
   959 => x"ffffff",
   960 => x"ffffff",
   961 => x"fff555",
   962 => x"555555",
   963 => x"555555",
   964 => x"555aaa",
   965 => x"ffffff",
   966 => x"ffffff",
   967 => x"ffffff",
   968 => x"ffffff",
   969 => x"ffffff",
   970 => x"ffffff",
   971 => x"ffffff",
   972 => x"ffffff",
   973 => x"ffffff",
   974 => x"ffffff",
   975 => x"ffffff",
   976 => x"ffffff",
   977 => x"ffffff",
   978 => x"ffffff",
   979 => x"ffffff",
   980 => x"ffffff",
   981 => x"ffffff",
   982 => x"ffffff",
   983 => x"ffffff",
   984 => x"ffffff",
   985 => x"ffffff",
   986 => x"ffffff",
   987 => x"ffffff",
   988 => x"ffffff",
   989 => x"ffffff",
   990 => x"ffffff",
   991 => x"ffffff",
   992 => x"ffffff",
   993 => x"ffffff",
   994 => x"ffffff",
   995 => x"ffffff",
   996 => x"ffffff",
   997 => x"ffffff",
   998 => x"ffffff",
   999 => x"ffffff",
   1000 => x"ffffff",
   1001 => x"ffffff",
   1002 => x"ffffff",
   1003 => x"ffffff",
   1004 => x"ffffff",
   1005 => x"ffffff",
   1006 => x"ffffff",
   1007 => x"ffffff",
   1008 => x"ffffff",
   1009 => x"ffffff",
   1010 => x"ffffff",
   1011 => x"ffffff",
   1012 => x"ffffff",
   1013 => x"ffffff",
   1014 => x"ffffff",
   1015 => x"ffffff",
   1016 => x"ffffff",
   1017 => x"ffffff",
   1018 => x"ffffff",
   1019 => x"ffffff",
   1020 => x"ffffff",
   1021 => x"ffffff",
   1022 => x"fffa95",
   1023 => x"000000",
   1024 => x"000000",
   1025 => x"000000",
   1026 => x"000000",
   1027 => x"015abf",
   1028 => x"ffffff",
   1029 => x"ffffff",
   1030 => x"ffffff",
   1031 => x"ffffff",
   1032 => x"ffffff",
   1033 => x"ffffff",
   1034 => x"ffffff",
   1035 => x"ffffff",
   1036 => x"ffffff",
   1037 => x"ffffff",
   1038 => x"ffffff",
   1039 => x"ffffff",
   1040 => x"ffffff",
   1041 => x"ffffff",
   1042 => x"ffffff",
   1043 => x"ffffff",
   1044 => x"ffffff",
   1045 => x"ffffff",
   1046 => x"ffffff",
   1047 => x"ffffff",
   1048 => x"ffffff",
   1049 => x"ffffff",
   1050 => x"ffffff",
   1051 => x"ffffff",
   1052 => x"ffffff",
   1053 => x"ffffff",
   1054 => x"ffffff",
   1055 => x"ffffff",
   1056 => x"ffffff",
   1057 => x"ffffff",
   1058 => x"ffffff",
   1059 => x"ffffff",
   1060 => x"ffffff",
   1061 => x"ffffff",
   1062 => x"ffffff",
   1063 => x"ffffff",
   1064 => x"ffffff",
   1065 => x"ffffff",
   1066 => x"ffffff",
   1067 => x"ffffff",
   1068 => x"ffffff",
   1069 => x"ffffff",
   1070 => x"a95abf",
   1071 => x"ffffff",
   1072 => x"ffffff",
   1073 => x"ffffff",
   1074 => x"ffffff",
   1075 => x"ffffff",
   1076 => x"ffffff",
   1077 => x"ffffff",
   1078 => x"ffffff",
   1079 => x"ffffff",
   1080 => x"ffffff",
   1081 => x"ffffff",
   1082 => x"ffffff",
   1083 => x"ffffff",
   1084 => x"ffffff",
   1085 => x"ffffff",
   1086 => x"ffffff",
   1087 => x"ffffff",
   1088 => x"ffffff",
   1089 => x"ffffff",
   1090 => x"ffffff",
   1091 => x"ffffff",
   1092 => x"ffffff",
   1093 => x"ffffff",
   1094 => x"ffffff",
   1095 => x"ffffff",
   1096 => x"ffffff",
   1097 => x"ffffff",
   1098 => x"ffffff",
   1099 => x"ffffff",
   1100 => x"ffffff",
   1101 => x"ffffff",
   1102 => x"ffffff",
   1103 => x"ffffff",
   1104 => x"ffffff",
   1105 => x"ffffff",
   1106 => x"ffffff",
   1107 => x"ffffff",
   1108 => x"ffffff",
   1109 => x"ffffff",
   1110 => x"ffffff",
   1111 => x"ffffff",
   1112 => x"ffffff",
   1113 => x"ffffff",
   1114 => x"ffffff",
   1115 => x"ffffff",
   1116 => x"ffffff",
   1117 => x"ffffff",
   1118 => x"ffffff",
   1119 => x"ffffff",
   1120 => x"ffffff",
   1121 => x"fff540",
   1122 => x"000000",
   1123 => x"000000",
   1124 => x"000000",
   1125 => x"555abf",
   1126 => x"ffffff",
   1127 => x"ffffff",
   1128 => x"ffffff",
   1129 => x"ffffff",
   1130 => x"ffffff",
   1131 => x"ffffff",
   1132 => x"ffffff",
   1133 => x"ffffff",
   1134 => x"ffffff",
   1135 => x"ffffff",
   1136 => x"ffffff",
   1137 => x"ffffff",
   1138 => x"ffffff",
   1139 => x"ffffff",
   1140 => x"ffffff",
   1141 => x"ffffff",
   1142 => x"ffffff",
   1143 => x"ffffff",
   1144 => x"ffffff",
   1145 => x"ffffff",
   1146 => x"ffffff",
   1147 => x"ffffff",
   1148 => x"ffffff",
   1149 => x"ffffff",
   1150 => x"ffffff",
   1151 => x"ffffff",
   1152 => x"ffffff",
   1153 => x"ffffff",
   1154 => x"ffffff",
   1155 => x"ffffff",
   1156 => x"ffffff",
   1157 => x"ffffff",
   1158 => x"ffffff",
   1159 => x"ffffff",
   1160 => x"ffffff",
   1161 => x"ffffff",
   1162 => x"ffffff",
   1163 => x"ffffff",
   1164 => x"ffffff",
   1165 => x"ffffff",
   1166 => x"ffffff",
   1167 => x"ffffff",
   1168 => x"ffffff",
   1169 => x"ffffff",
   1170 => x"ffffff",
   1171 => x"ffffff",
   1172 => x"ffffff",
   1173 => x"ffffff",
   1174 => x"ffffff",
   1175 => x"ffffff",
   1176 => x"ffffff",
   1177 => x"ffffff",
   1178 => x"ffffff",
   1179 => x"ffffff",
   1180 => x"ffffff",
   1181 => x"ffffff",
   1182 => x"fea540",
   1183 => x"000000",
   1184 => x"555aaa",
   1185 => x"aaaa95",
   1186 => x"540000",
   1187 => x"00057f",
   1188 => x"ffffff",
   1189 => x"ffffff",
   1190 => x"ffffff",
   1191 => x"ffffff",
   1192 => x"ffffff",
   1193 => x"ffffff",
   1194 => x"ffffff",
   1195 => x"ffffff",
   1196 => x"ffffff",
   1197 => x"ffffff",
   1198 => x"ffffff",
   1199 => x"ffffff",
   1200 => x"ffffff",
   1201 => x"ffffff",
   1202 => x"ffffff",
   1203 => x"ffffff",
   1204 => x"ffffff",
   1205 => x"ffffff",
   1206 => x"ffffff",
   1207 => x"ffffff",
   1208 => x"ffffff",
   1209 => x"ffffff",
   1210 => x"ffffff",
   1211 => x"ffffff",
   1212 => x"ffffff",
   1213 => x"ffffff",
   1214 => x"ffffff",
   1215 => x"ffffff",
   1216 => x"ffffff",
   1217 => x"ffffff",
   1218 => x"ffffff",
   1219 => x"ffffff",
   1220 => x"ffffff",
   1221 => x"ffffff",
   1222 => x"ffffff",
   1223 => x"ffffff",
   1224 => x"ffffff",
   1225 => x"ffffff",
   1226 => x"ffffff",
   1227 => x"ffffff",
   1228 => x"ffffff",
   1229 => x"ffffea",
   1230 => x"56afff",
   1231 => x"ffffff",
   1232 => x"ffffff",
   1233 => x"ffffff",
   1234 => x"ffffff",
   1235 => x"ffffff",
   1236 => x"ffffff",
   1237 => x"ffffff",
   1238 => x"ffffff",
   1239 => x"ffffff",
   1240 => x"ffffff",
   1241 => x"ffffff",
   1242 => x"ffffff",
   1243 => x"ffffff",
   1244 => x"ffffff",
   1245 => x"ffffff",
   1246 => x"ffffff",
   1247 => x"ffffff",
   1248 => x"ffffff",
   1249 => x"ffffff",
   1250 => x"ffffff",
   1251 => x"ffffff",
   1252 => x"ffffff",
   1253 => x"ffffff",
   1254 => x"ffffff",
   1255 => x"ffffff",
   1256 => x"ffffff",
   1257 => x"ffffff",
   1258 => x"ffffff",
   1259 => x"ffffff",
   1260 => x"ffffff",
   1261 => x"ffffff",
   1262 => x"ffffff",
   1263 => x"ffffff",
   1264 => x"ffffff",
   1265 => x"ffffff",
   1266 => x"ffffff",
   1267 => x"ffffff",
   1268 => x"ffffff",
   1269 => x"ffffff",
   1270 => x"ffffff",
   1271 => x"ffffff",
   1272 => x"ffffff",
   1273 => x"ffffff",
   1274 => x"ffffff",
   1275 => x"ffffff",
   1276 => x"ffffff",
   1277 => x"ffffff",
   1278 => x"ffffff",
   1279 => x"ffffff",
   1280 => x"ffffff",
   1281 => x"fff540",
   1282 => x"000000",
   1283 => x"000000",
   1284 => x"000000",
   1285 => x"00056a",
   1286 => x"ffffff",
   1287 => x"ffffff",
   1288 => x"ffffff",
   1289 => x"ffffff",
   1290 => x"ffffff",
   1291 => x"ffffff",
   1292 => x"ffffff",
   1293 => x"ffffff",
   1294 => x"ffffff",
   1295 => x"ffffff",
   1296 => x"ffffff",
   1297 => x"ffffff",
   1298 => x"ffffff",
   1299 => x"ffffff",
   1300 => x"ffffff",
   1301 => x"ffffff",
   1302 => x"ffffff",
   1303 => x"ffffff",
   1304 => x"ffffff",
   1305 => x"ffffff",
   1306 => x"ffffff",
   1307 => x"ffffff",
   1308 => x"ffffff",
   1309 => x"ffffff",
   1310 => x"ffffff",
   1311 => x"ffffff",
   1312 => x"ffffff",
   1313 => x"ffffff",
   1314 => x"ffffff",
   1315 => x"ffffff",
   1316 => x"ffffff",
   1317 => x"ffffff",
   1318 => x"ffffff",
   1319 => x"ffffff",
   1320 => x"ffffff",
   1321 => x"ffffff",
   1322 => x"ffffff",
   1323 => x"ffffff",
   1324 => x"ffffff",
   1325 => x"ffffff",
   1326 => x"ffffff",
   1327 => x"ffffff",
   1328 => x"ffffff",
   1329 => x"ffffff",
   1330 => x"ffffff",
   1331 => x"ffffff",
   1332 => x"ffffff",
   1333 => x"ffffff",
   1334 => x"ffffff",
   1335 => x"ffffff",
   1336 => x"ffffff",
   1337 => x"ffffff",
   1338 => x"ffffff",
   1339 => x"ffffff",
   1340 => x"ffffff",
   1341 => x"ffffff",
   1342 => x"a95000",
   1343 => x"00056a",
   1344 => x"abffff",
   1345 => x"ffffff",
   1346 => x"feaa95",
   1347 => x"00003f",
   1348 => x"ffffff",
   1349 => x"ffffff",
   1350 => x"ffffff",
   1351 => x"ffffff",
   1352 => x"ffffff",
   1353 => x"ffffff",
   1354 => x"ffffff",
   1355 => x"ffffff",
   1356 => x"ffffff",
   1357 => x"ffffff",
   1358 => x"ffffff",
   1359 => x"ffffff",
   1360 => x"ffffff",
   1361 => x"ffffff",
   1362 => x"ffffff",
   1363 => x"ffffff",
   1364 => x"ffffff",
   1365 => x"ffffff",
   1366 => x"ffffff",
   1367 => x"ffffff",
   1368 => x"ffffff",
   1369 => x"ffffff",
   1370 => x"ffffff",
   1371 => x"ffffff",
   1372 => x"ffffff",
   1373 => x"ffffff",
   1374 => x"ffffff",
   1375 => x"ffffff",
   1376 => x"ffffff",
   1377 => x"ffffff",
   1378 => x"ffffff",
   1379 => x"ffffff",
   1380 => x"ffffff",
   1381 => x"ffffff",
   1382 => x"ffffff",
   1383 => x"ffffff",
   1384 => x"ffffff",
   1385 => x"ffffff",
   1386 => x"ffffff",
   1387 => x"ffffff",
   1388 => x"ffffff",
   1389 => x"fffa95",
   1390 => x"abffff",
   1391 => x"ffffff",
   1392 => x"ffffff",
   1393 => x"ffffff",
   1394 => x"ffffff",
   1395 => x"ffffff",
   1396 => x"ffffff",
   1397 => x"ffffff",
   1398 => x"ffffff",
   1399 => x"ffffff",
   1400 => x"ffffff",
   1401 => x"ffffff",
   1402 => x"ffffff",
   1403 => x"ffffff",
   1404 => x"ffffff",
   1405 => x"ffffff",
   1406 => x"ffffff",
   1407 => x"ffffff",
   1408 => x"ffffff",
   1409 => x"ffffff",
   1410 => x"ffffff",
   1411 => x"ffffff",
   1412 => x"ffffff",
   1413 => x"ffffff",
   1414 => x"ffffff",
   1415 => x"ffffff",
   1416 => x"ffffff",
   1417 => x"ffffff",
   1418 => x"ffffff",
   1419 => x"ffffff",
   1420 => x"ffffff",
   1421 => x"ffffff",
   1422 => x"ffffff",
   1423 => x"ffffff",
   1424 => x"ffffff",
   1425 => x"ffffff",
   1426 => x"ffffff",
   1427 => x"ffffff",
   1428 => x"ffffff",
   1429 => x"ffffff",
   1430 => x"ffffff",
   1431 => x"ffffff",
   1432 => x"ffffff",
   1433 => x"ffffff",
   1434 => x"ffffff",
   1435 => x"ffffff",
   1436 => x"ffffff",
   1437 => x"ffffff",
   1438 => x"ffffff",
   1439 => x"ffffff",
   1440 => x"ffffff",
   1441 => x"fff540",
   1442 => x"000555",
   1443 => x"555555",
   1444 => x"555000",
   1445 => x"000015",
   1446 => x"abffff",
   1447 => x"ffffff",
   1448 => x"ffffff",
   1449 => x"ffffff",
   1450 => x"ffffff",
   1451 => x"ffffff",
   1452 => x"ffffff",
   1453 => x"ffffff",
   1454 => x"ffffff",
   1455 => x"ffffff",
   1456 => x"ffffff",
   1457 => x"ffffff",
   1458 => x"ffffff",
   1459 => x"ffffff",
   1460 => x"ffffff",
   1461 => x"ffffff",
   1462 => x"ffffff",
   1463 => x"ffffff",
   1464 => x"ffffff",
   1465 => x"ffffff",
   1466 => x"ffffff",
   1467 => x"ffffff",
   1468 => x"ffffff",
   1469 => x"ffffff",
   1470 => x"ffffff",
   1471 => x"ffffff",
   1472 => x"ffffff",
   1473 => x"ffffff",
   1474 => x"ffffff",
   1475 => x"ffffff",
   1476 => x"ffffff",
   1477 => x"ffffff",
   1478 => x"ffffff",
   1479 => x"ffffff",
   1480 => x"ffffff",
   1481 => x"ffffff",
   1482 => x"ffffff",
   1483 => x"ffffff",
   1484 => x"ffffff",
   1485 => x"ffffff",
   1486 => x"ffffff",
   1487 => x"ffffff",
   1488 => x"ffffff",
   1489 => x"ffffff",
   1490 => x"ffffff",
   1491 => x"ffffff",
   1492 => x"ffffff",
   1493 => x"ffffff",
   1494 => x"ffffff",
   1495 => x"ffffff",
   1496 => x"ffffff",
   1497 => x"ffffff",
   1498 => x"ffffff",
   1499 => x"ffffff",
   1500 => x"ffffff",
   1501 => x"ffffff",
   1502 => x"540000",
   1503 => x"02afff",
   1504 => x"ffffff",
   1505 => x"ffffff",
   1506 => x"ffffea",
   1507 => x"a8003f",
   1508 => x"ffffff",
   1509 => x"ffffff",
   1510 => x"ffffff",
   1511 => x"ffffff",
   1512 => x"ffffff",
   1513 => x"ffffff",
   1514 => x"ffffff",
   1515 => x"ffffff",
   1516 => x"ffffff",
   1517 => x"ffffff",
   1518 => x"ffffff",
   1519 => x"ffffff",
   1520 => x"ffffff",
   1521 => x"ffffff",
   1522 => x"ffffff",
   1523 => x"ffffff",
   1524 => x"ffffff",
   1525 => x"ffffff",
   1526 => x"ffffff",
   1527 => x"ffffff",
   1528 => x"ffffff",
   1529 => x"ffffff",
   1530 => x"ffffff",
   1531 => x"ffffff",
   1532 => x"ffffff",
   1533 => x"ffffff",
   1534 => x"ffffff",
   1535 => x"ffffff",
   1536 => x"ffffff",
   1537 => x"ffffff",
   1538 => x"ffffff",
   1539 => x"ffffff",
   1540 => x"ffffff",
   1541 => x"ffffff",
   1542 => x"ffffff",
   1543 => x"ffffff",
   1544 => x"ffffff",
   1545 => x"ffffff",
   1546 => x"ffffff",
   1547 => x"ffffff",
   1548 => x"ffffff",
   1549 => x"fea56a",
   1550 => x"ffffff",
   1551 => x"ffffff",
   1552 => x"ffffff",
   1553 => x"ffffff",
   1554 => x"ffffff",
   1555 => x"ffffff",
   1556 => x"ffffff",
   1557 => x"ffffff",
   1558 => x"ffffff",
   1559 => x"ffffff",
   1560 => x"ffffff",
   1561 => x"ffffff",
   1562 => x"ffffff",
   1563 => x"ffffff",
   1564 => x"ffffff",
   1565 => x"ffffff",
   1566 => x"ffffff",
   1567 => x"ffffff",
   1568 => x"ffffff",
   1569 => x"ffffff",
   1570 => x"ffffff",
   1571 => x"ffffff",
   1572 => x"ffffff",
   1573 => x"ffffff",
   1574 => x"ffffff",
   1575 => x"ffffff",
   1576 => x"ffffff",
   1577 => x"ffffff",
   1578 => x"ffffff",
   1579 => x"ffffff",
   1580 => x"ffffff",
   1581 => x"ffffff",
   1582 => x"ffffff",
   1583 => x"ffffff",
   1584 => x"ffffff",
   1585 => x"ffffff",
   1586 => x"ffffff",
   1587 => x"ffffff",
   1588 => x"ffffff",
   1589 => x"ffffff",
   1590 => x"ffffff",
   1591 => x"ffffff",
   1592 => x"ffffff",
   1593 => x"ffffff",
   1594 => x"ffffff",
   1595 => x"ffffff",
   1596 => x"ffffff",
   1597 => x"ffffff",
   1598 => x"ffffff",
   1599 => x"ffffff",
   1600 => x"ffffff",
   1601 => x"fff540",
   1602 => x"000abf",
   1603 => x"ffffff",
   1604 => x"feaa95",
   1605 => x"000000",
   1606 => x"57ffff",
   1607 => x"ffffff",
   1608 => x"ffffff",
   1609 => x"ffffff",
   1610 => x"ffffff",
   1611 => x"ffffff",
   1612 => x"ffffff",
   1613 => x"ffffff",
   1614 => x"ffffff",
   1615 => x"ffffff",
   1616 => x"ffffff",
   1617 => x"ffffff",
   1618 => x"ffffff",
   1619 => x"ffffff",
   1620 => x"ffffff",
   1621 => x"ffffff",
   1622 => x"ffffff",
   1623 => x"ffffff",
   1624 => x"ffffff",
   1625 => x"ffffff",
   1626 => x"ffffff",
   1627 => x"ffffff",
   1628 => x"ffffff",
   1629 => x"ffffff",
   1630 => x"ffffff",
   1631 => x"ffffff",
   1632 => x"ffffff",
   1633 => x"ffffff",
   1634 => x"ffffff",
   1635 => x"ffffff",
   1636 => x"ffffff",
   1637 => x"ffffff",
   1638 => x"ffffff",
   1639 => x"ffffff",
   1640 => x"ffffff",
   1641 => x"ffffff",
   1642 => x"ffffff",
   1643 => x"ffffff",
   1644 => x"ffffff",
   1645 => x"ffffff",
   1646 => x"ffffff",
   1647 => x"ffffff",
   1648 => x"ffffff",
   1649 => x"ffffff",
   1650 => x"ffffff",
   1651 => x"ffffff",
   1652 => x"ffffff",
   1653 => x"ffffff",
   1654 => x"ffffff",
   1655 => x"ffffff",
   1656 => x"ffffff",
   1657 => x"ffffff",
   1658 => x"ffffff",
   1659 => x"ffffff",
   1660 => x"ffffff",
   1661 => x"ffffd5",
   1662 => x"000000",
   1663 => x"abffff",
   1664 => x"ffffff",
   1665 => x"ffffff",
   1666 => x"ffffff",
   1667 => x"fea57f",
   1668 => x"ffffff",
   1669 => x"ffffff",
   1670 => x"ffffff",
   1671 => x"ffffff",
   1672 => x"ffffff",
   1673 => x"ffffff",
   1674 => x"ffffff",
   1675 => x"ffffff",
   1676 => x"ffffff",
   1677 => x"ffffff",
   1678 => x"ffffff",
   1679 => x"ffffff",
   1680 => x"ffffff",
   1681 => x"ffffff",
   1682 => x"ffffff",
   1683 => x"ffffff",
   1684 => x"ffffff",
   1685 => x"ffffff",
   1686 => x"ffffff",
   1687 => x"ffffff",
   1688 => x"ffffff",
   1689 => x"ffffff",
   1690 => x"ffffff",
   1691 => x"ffffff",
   1692 => x"ffffff",
   1693 => x"ffffff",
   1694 => x"ffffff",
   1695 => x"ffffff",
   1696 => x"ffffff",
   1697 => x"ffffff",
   1698 => x"ffffff",
   1699 => x"ffffff",
   1700 => x"ffffff",
   1701 => x"ffffff",
   1702 => x"ffffff",
   1703 => x"ffffff",
   1704 => x"ffffff",
   1705 => x"ffffff",
   1706 => x"ffffff",
   1707 => x"ffffff",
   1708 => x"ffffff",
   1709 => x"a95abf",
   1710 => x"ffffff",
   1711 => x"ffffff",
   1712 => x"ffffff",
   1713 => x"ffffff",
   1714 => x"ffffff",
   1715 => x"ffffff",
   1716 => x"ffffff",
   1717 => x"ffffff",
   1718 => x"ffffff",
   1719 => x"ffffff",
   1720 => x"ffffff",
   1721 => x"ffffff",
   1722 => x"ffffff",
   1723 => x"ffffff",
   1724 => x"ffffff",
   1725 => x"ffffff",
   1726 => x"ffffff",
   1727 => x"ffffff",
   1728 => x"ffffff",
   1729 => x"ffffff",
   1730 => x"ffffff",
   1731 => x"ffffff",
   1732 => x"ffffff",
   1733 => x"ffffff",
   1734 => x"ffffff",
   1735 => x"ffffff",
   1736 => x"ffffff",
   1737 => x"ffffff",
   1738 => x"ffffff",
   1739 => x"ffffff",
   1740 => x"ffffff",
   1741 => x"ffffff",
   1742 => x"ffffff",
   1743 => x"ffffff",
   1744 => x"ffffff",
   1745 => x"ffffff",
   1746 => x"ffffff",
   1747 => x"ffffff",
   1748 => x"ffffff",
   1749 => x"ffffff",
   1750 => x"ffffff",
   1751 => x"ffffff",
   1752 => x"ffffff",
   1753 => x"ffffff",
   1754 => x"ffffff",
   1755 => x"ffffff",
   1756 => x"ffffff",
   1757 => x"ffffff",
   1758 => x"ffffff",
   1759 => x"ffffff",
   1760 => x"ffffff",
   1761 => x"fff540",
   1762 => x"000abf",
   1763 => x"ffffff",
   1764 => x"ffffea",
   1765 => x"540000",
   1766 => x"02afff",
   1767 => x"ffffff",
   1768 => x"ffffff",
   1769 => x"ffffff",
   1770 => x"ffffff",
   1771 => x"ffffff",
   1772 => x"ffffff",
   1773 => x"ffffff",
   1774 => x"ffffff",
   1775 => x"ffffff",
   1776 => x"ffffff",
   1777 => x"ffffff",
   1778 => x"ffffff",
   1779 => x"ffffff",
   1780 => x"ffffff",
   1781 => x"ffffff",
   1782 => x"ffffff",
   1783 => x"ffffff",
   1784 => x"ffffff",
   1785 => x"ffffff",
   1786 => x"ffffff",
   1787 => x"ffffff",
   1788 => x"ffffff",
   1789 => x"ffffff",
   1790 => x"ffffff",
   1791 => x"ffffff",
   1792 => x"ffffff",
   1793 => x"ffffff",
   1794 => x"ffffff",
   1795 => x"ffffff",
   1796 => x"ffffff",
   1797 => x"ffffff",
   1798 => x"ffffff",
   1799 => x"ffffff",
   1800 => x"ffffff",
   1801 => x"ffffff",
   1802 => x"ffffff",
   1803 => x"ffffff",
   1804 => x"ffffff",
   1805 => x"ffffff",
   1806 => x"ffffff",
   1807 => x"ffffff",
   1808 => x"ffffff",
   1809 => x"ffffff",
   1810 => x"ffffff",
   1811 => x"ffffff",
   1812 => x"ffffff",
   1813 => x"ffffff",
   1814 => x"ffffff",
   1815 => x"ffffff",
   1816 => x"ffffff",
   1817 => x"ffffff",
   1818 => x"ffffff",
   1819 => x"ffffff",
   1820 => x"ffffff",
   1821 => x"ffffd5",
   1822 => x"000015",
   1823 => x"ffffff",
   1824 => x"ffffff",
   1825 => x"ffffff",
   1826 => x"ffffff",
   1827 => x"ffffff",
   1828 => x"ffffff",
   1829 => x"ffffff",
   1830 => x"ffffff",
   1831 => x"ffffff",
   1832 => x"ffffff",
   1833 => x"ffffff",
   1834 => x"ffffff",
   1835 => x"ffffff",
   1836 => x"ffffff",
   1837 => x"ffffff",
   1838 => x"ffffff",
   1839 => x"ffffff",
   1840 => x"ffffff",
   1841 => x"ffffff",
   1842 => x"ffffff",
   1843 => x"ffffff",
   1844 => x"ffffff",
   1845 => x"ffffff",
   1846 => x"ffffff",
   1847 => x"ffffff",
   1848 => x"ffffff",
   1849 => x"ffffff",
   1850 => x"ffffff",
   1851 => x"ffffff",
   1852 => x"ffffff",
   1853 => x"ffffff",
   1854 => x"ffffff",
   1855 => x"ffffff",
   1856 => x"ffffff",
   1857 => x"ffffff",
   1858 => x"ffffff",
   1859 => x"ffffff",
   1860 => x"ffffff",
   1861 => x"ffffff",
   1862 => x"ffffff",
   1863 => x"ffffff",
   1864 => x"ffffff",
   1865 => x"ffffff",
   1866 => x"ffffff",
   1867 => x"ffffff",
   1868 => x"ffffea",
   1869 => x"56afff",
   1870 => x"ffffff",
   1871 => x"ffffff",
   1872 => x"ffffff",
   1873 => x"ffffff",
   1874 => x"ffffff",
   1875 => x"ffffff",
   1876 => x"ffffff",
   1877 => x"ffffff",
   1878 => x"ffffff",
   1879 => x"ffffff",
   1880 => x"ffffff",
   1881 => x"ffffff",
   1882 => x"ffffff",
   1883 => x"ffffff",
   1884 => x"ffffff",
   1885 => x"ffffff",
   1886 => x"ffffff",
   1887 => x"ffffff",
   1888 => x"ffffff",
   1889 => x"ffffff",
   1890 => x"ffffff",
   1891 => x"ffffff",
   1892 => x"ffffff",
   1893 => x"ffffff",
   1894 => x"ffffff",
   1895 => x"ffffff",
   1896 => x"ffffff",
   1897 => x"ffffff",
   1898 => x"ffffff",
   1899 => x"ffffff",
   1900 => x"ffffff",
   1901 => x"ffffff",
   1902 => x"ffffff",
   1903 => x"ffffff",
   1904 => x"ffffff",
   1905 => x"ffffff",
   1906 => x"ffffff",
   1907 => x"ffffff",
   1908 => x"ffffff",
   1909 => x"ffffff",
   1910 => x"ffffff",
   1911 => x"ffffff",
   1912 => x"ffffff",
   1913 => x"ffffff",
   1914 => x"ffffff",
   1915 => x"ffffff",
   1916 => x"ffffff",
   1917 => x"ffffff",
   1918 => x"ffffff",
   1919 => x"ffffff",
   1920 => x"ffffff",
   1921 => x"fff540",
   1922 => x"000abf",
   1923 => x"ffffff",
   1924 => x"ffffff",
   1925 => x"a80000",
   1926 => x"02afff",
   1927 => x"ffffff",
   1928 => x"ffffff",
   1929 => x"ffffff",
   1930 => x"ffffff",
   1931 => x"ffffff",
   1932 => x"ffffff",
   1933 => x"ffffff",
   1934 => x"ffffff",
   1935 => x"ffffff",
   1936 => x"ffffff",
   1937 => x"ffffff",
   1938 => x"ffffff",
   1939 => x"ffffff",
   1940 => x"ffaeba",
   1941 => x"eb5d75",
   1942 => x"d75d75",
   1943 => x"d75d75",
   1944 => x"d75d75",
   1945 => x"d75eba",
   1946 => x"ebaebf",
   1947 => x"ffffff",
   1948 => x"ffffff",
   1949 => x"ffffff",
   1950 => x"ffffff",
   1951 => x"ffffff",
   1952 => x"ffffff",
   1953 => x"ffffff",
   1954 => x"ffffff",
   1955 => x"ffffff",
   1956 => x"ffffff",
   1957 => x"ffffff",
   1958 => x"ffffff",
   1959 => x"ffffff",
   1960 => x"ffffff",
   1961 => x"ffffff",
   1962 => x"baebae",
   1963 => x"75d75d",
   1964 => x"75d75d",
   1965 => x"75d75d",
   1966 => x"75d75d",
   1967 => x"76ebae",
   1968 => x"baefff",
   1969 => x"ffffff",
   1970 => x"ffffff",
   1971 => x"ffffff",
   1972 => x"ffffff",
   1973 => x"ffffff",
   1974 => x"ffffff",
   1975 => x"ffffff",
   1976 => x"ffffff",
   1977 => x"ffffff",
   1978 => x"ffffff",
   1979 => x"ffffff",
   1980 => x"ffffff",
   1981 => x"fffa80",
   1982 => x"00056a",
   1983 => x"ffffff",
   1984 => x"ffffff",
   1985 => x"ffffff",
   1986 => x"ffffff",
   1987 => x"ffffff",
   1988 => x"ffffff",
   1989 => x"ffffff",
   1990 => x"ffffff",
   1991 => x"ffffff",
   1992 => x"ffffff",
   1993 => x"ffffff",
   1994 => x"ffffff",
   1995 => x"ffffff",
   1996 => x"ffffff",
   1997 => x"ffffff",
   1998 => x"ffffff",
   1999 => x"ffffff",
   2000 => x"ffffff",
   2001 => x"ffffff",
   2002 => x"ffffff",
   2003 => x"ffffff",
   2004 => x"ffffff",
   2005 => x"ffffff",
   2006 => x"ffffff",
   2007 => x"ffffff",
   2008 => x"ffffff",
   2009 => x"ffffff",
   2010 => x"ffffff",
   2011 => x"ffffff",
   2012 => x"ffffff",
   2013 => x"ffffff",
   2014 => x"ffffff",
   2015 => x"ffffff",
   2016 => x"ffffff",
   2017 => x"ffffff",
   2018 => x"ffffff",
   2019 => x"ffffff",
   2020 => x"ffffff",
   2021 => x"ffffff",
   2022 => x"ffffff",
   2023 => x"ffffff",
   2024 => x"ffffff",
   2025 => x"ffffff",
   2026 => x"ffffff",
   2027 => x"ffffff",
   2028 => x"fffa95",
   2029 => x"abffff",
   2030 => x"ffffff",
   2031 => x"ffffff",
   2032 => x"ffffff",
   2033 => x"ffffff",
   2034 => x"ffffff",
   2035 => x"ffffff",
   2036 => x"ffffff",
   2037 => x"ffffff",
   2038 => x"ffffff",
   2039 => x"ffffff",
   2040 => x"ffffff",
   2041 => x"ffffff",
   2042 => x"ffffff",
   2043 => x"ffffff",
   2044 => x"ffffff",
   2045 => x"ffffff",
   2046 => x"ffffff",
   2047 => x"ffffff",
   2048 => x"ffffff",
   2049 => x"ffffff",
   2050 => x"ffffff",
   2051 => x"ffffff",
   2052 => x"ffffff",
   2053 => x"ffffff",
   2054 => x"ffffff",
   2055 => x"ffffff",
   2056 => x"ffffff",
   2057 => x"ffffff",
   2058 => x"ffffff",
   2059 => x"ffffff",
   2060 => x"ffffff",
   2061 => x"ffffff",
   2062 => x"ffffff",
   2063 => x"ffffff",
   2064 => x"ffffff",
   2065 => x"ffffff",
   2066 => x"ffffff",
   2067 => x"ffffff",
   2068 => x"ffffff",
   2069 => x"ffffff",
   2070 => x"ffffff",
   2071 => x"ffffff",
   2072 => x"ffffff",
   2073 => x"ffffff",
   2074 => x"ffffff",
   2075 => x"ffffff",
   2076 => x"ffffff",
   2077 => x"ffffff",
   2078 => x"ffffff",
   2079 => x"ffffff",
   2080 => x"ffffff",
   2081 => x"fff540",
   2082 => x"000abf",
   2083 => x"ffffff",
   2084 => x"ffffff",
   2085 => x"fd5000",
   2086 => x"015fff",
   2087 => x"ffffff",
   2088 => x"ffffff",
   2089 => x"ffffff",
   2090 => x"ffffff",
   2091 => x"ffffff",
   2092 => x"ffffff",
   2093 => x"ffffff",
   2094 => x"ffffff",
   2095 => x"ffffff",
   2096 => x"ffffff",
   2097 => x"ffffff",
   2098 => x"fffffa",
   2099 => x"ebad75",
   2100 => x"d75c30",
   2101 => x"c30c30",
   2102 => x"c30c30",
   2103 => x"c30c30",
   2104 => x"c30c30",
   2105 => x"c30c30",
   2106 => x"c35d75",
   2107 => x"d7aeba",
   2108 => x"ebffff",
   2109 => x"ffffff",
   2110 => x"ffffff",
   2111 => x"ffffff",
   2112 => x"ffffff",
   2113 => x"ffffff",
   2114 => x"ffffff",
   2115 => x"ffffff",
   2116 => x"ffffff",
   2117 => x"ffffff",
   2118 => x"ffffff",
   2119 => x"ffffff",
   2120 => x"fffbae",
   2121 => x"bae75d",
   2122 => x"75d30c",
   2123 => x"30c30c",
   2124 => x"30c30c",
   2125 => x"30c30c",
   2126 => x"30c30c",
   2127 => x"30c30c",
   2128 => x"75d75d",
   2129 => x"baebae",
   2130 => x"ffffff",
   2131 => x"ffffff",
   2132 => x"ffffff",
   2133 => x"ffffff",
   2134 => x"ffffff",
   2135 => x"ffffff",
   2136 => x"ffffff",
   2137 => x"ffffff",
   2138 => x"ffffff",
   2139 => x"ffffff",
   2140 => x"ffffff",
   2141 => x"fff540",
   2142 => x"00057f",
   2143 => x"ffffff",
   2144 => x"ffffff",
   2145 => x"ffffff",
   2146 => x"ffffff",
   2147 => x"ffffff",
   2148 => x"ffffff",
   2149 => x"ffffff",
   2150 => x"ffffff",
   2151 => x"ffffff",
   2152 => x"ffffff",
   2153 => x"ffffff",
   2154 => x"ffffff",
   2155 => x"ffffff",
   2156 => x"ffffff",
   2157 => x"ffffff",
   2158 => x"ffffff",
   2159 => x"ffffff",
   2160 => x"ffffff",
   2161 => x"ffffff",
   2162 => x"ffffff",
   2163 => x"ffffff",
   2164 => x"ffffff",
   2165 => x"ffffff",
   2166 => x"ffffff",
   2167 => x"ffffff",
   2168 => x"ffffff",
   2169 => x"ffffff",
   2170 => x"ffffff",
   2171 => x"ffffff",
   2172 => x"ffffff",
   2173 => x"ffffff",
   2174 => x"ffffff",
   2175 => x"ffffff",
   2176 => x"ffffff",
   2177 => x"ffffff",
   2178 => x"ffffff",
   2179 => x"ffffff",
   2180 => x"ffffff",
   2181 => x"ffffff",
   2182 => x"ffffff",
   2183 => x"ffffff",
   2184 => x"ffffff",
   2185 => x"ffffff",
   2186 => x"ffffff",
   2187 => x"ffffff",
   2188 => x"fea56a",
   2189 => x"ffffff",
   2190 => x"ffffff",
   2191 => x"ffffff",
   2192 => x"ffffff",
   2193 => x"ffffff",
   2194 => x"ffffff",
   2195 => x"ffffff",
   2196 => x"ffffff",
   2197 => x"ffffff",
   2198 => x"ffffff",
   2199 => x"ffffff",
   2200 => x"ffffff",
   2201 => x"ffffff",
   2202 => x"ffffff",
   2203 => x"ffffff",
   2204 => x"ffffff",
   2205 => x"ffffff",
   2206 => x"ffffff",
   2207 => x"ffffff",
   2208 => x"ffffff",
   2209 => x"ffffff",
   2210 => x"ffffff",
   2211 => x"ffffff",
   2212 => x"ffffff",
   2213 => x"ffffff",
   2214 => x"ffffff",
   2215 => x"ffffff",
   2216 => x"ffffff",
   2217 => x"ffffff",
   2218 => x"ffffff",
   2219 => x"ffffff",
   2220 => x"ffffff",
   2221 => x"ffffff",
   2222 => x"ffffff",
   2223 => x"ffffff",
   2224 => x"ffffff",
   2225 => x"ffffff",
   2226 => x"ffffff",
   2227 => x"ffffff",
   2228 => x"ffffff",
   2229 => x"ffffff",
   2230 => x"ffffff",
   2231 => x"ffffff",
   2232 => x"ffffff",
   2233 => x"ffffff",
   2234 => x"ffffff",
   2235 => x"ffffff",
   2236 => x"ffffff",
   2237 => x"ffffff",
   2238 => x"ffffff",
   2239 => x"ffffff",
   2240 => x"ffffff",
   2241 => x"fff540",
   2242 => x"000abf",
   2243 => x"ffffff",
   2244 => x"ffffff",
   2245 => x"fd5000",
   2246 => x"015fff",
   2247 => x"ffffff",
   2248 => x"ffffff",
   2249 => x"ffffff",
   2250 => x"ffffff",
   2251 => x"ffffff",
   2252 => x"ffffff",
   2253 => x"ffffff",
   2254 => x"ffffff",
   2255 => x"ffffff",
   2256 => x"ffffff",
   2257 => x"fffffa",
   2258 => x"eb5d75",
   2259 => x"c30c30",
   2260 => x"c30c30",
   2261 => x"c30c30",
   2262 => x"c30c30",
   2263 => x"c30c30",
   2264 => x"c30c30",
   2265 => x"c30c30",
   2266 => x"c30c30",
   2267 => x"c30c35",
   2268 => x"d75eba",
   2269 => x"ebffff",
   2270 => x"ffffff",
   2271 => x"ffffff",
   2272 => x"ffffff",
   2273 => x"ffffff",
   2274 => x"ffffff",
   2275 => x"ffffff",
   2276 => x"ffffff",
   2277 => x"ffffff",
   2278 => x"ffffff",
   2279 => x"fffbae",
   2280 => x"75d74c",
   2281 => x"30c30c",
   2282 => x"30c30c",
   2283 => x"30c30c",
   2284 => x"30c30c",
   2285 => x"30c30c",
   2286 => x"30c30c",
   2287 => x"30c30c",
   2288 => x"30c30c",
   2289 => x"30c31d",
   2290 => x"76ebae",
   2291 => x"ffffff",
   2292 => x"ffffff",
   2293 => x"ffffff",
   2294 => x"ffffff",
   2295 => x"ffffff",
   2296 => x"ffffff",
   2297 => x"ffffff",
   2298 => x"ffffff",
   2299 => x"ffffff",
   2300 => x"ffffff",
   2301 => x"fea540",
   2302 => x"000abf",
   2303 => x"ffffff",
   2304 => x"ffffff",
   2305 => x"ffffff",
   2306 => x"ffffff",
   2307 => x"ffffff",
   2308 => x"ffffff",
   2309 => x"ffffff",
   2310 => x"ffffff",
   2311 => x"ffffff",
   2312 => x"ffffff",
   2313 => x"ffffff",
   2314 => x"ffffff",
   2315 => x"ffffff",
   2316 => x"ffffff",
   2317 => x"ffffff",
   2318 => x"ffffff",
   2319 => x"ffffff",
   2320 => x"ffffff",
   2321 => x"ffffff",
   2322 => x"ffffff",
   2323 => x"ffffff",
   2324 => x"ffffff",
   2325 => x"ffffff",
   2326 => x"ffffff",
   2327 => x"ffffff",
   2328 => x"ffffff",
   2329 => x"ffffff",
   2330 => x"ffffff",
   2331 => x"ffffff",
   2332 => x"ffffff",
   2333 => x"ffffff",
   2334 => x"ffffff",
   2335 => x"ffffff",
   2336 => x"ffffff",
   2337 => x"ffffff",
   2338 => x"ffffff",
   2339 => x"ffffff",
   2340 => x"ffffff",
   2341 => x"ffffff",
   2342 => x"ffffff",
   2343 => x"ffffff",
   2344 => x"ffffff",
   2345 => x"ffffff",
   2346 => x"ffffff",
   2347 => x"ffffff",
   2348 => x"a95abf",
   2349 => x"ffffff",
   2350 => x"ffffff",
   2351 => x"ffffff",
   2352 => x"ffffff",
   2353 => x"ffffff",
   2354 => x"ffffff",
   2355 => x"ffffff",
   2356 => x"ffffff",
   2357 => x"ffffff",
   2358 => x"ffffff",
   2359 => x"ffffff",
   2360 => x"ffffff",
   2361 => x"ffffff",
   2362 => x"ffffff",
   2363 => x"ffffff",
   2364 => x"ffffff",
   2365 => x"ffffff",
   2366 => x"ffffff",
   2367 => x"ffffff",
   2368 => x"ffffff",
   2369 => x"ffffff",
   2370 => x"ffffff",
   2371 => x"ffffff",
   2372 => x"ffffff",
   2373 => x"ffffff",
   2374 => x"ffffff",
   2375 => x"ffffff",
   2376 => x"ffffff",
   2377 => x"ffffff",
   2378 => x"ffffff",
   2379 => x"ffffff",
   2380 => x"ffffff",
   2381 => x"ffffff",
   2382 => x"ffffff",
   2383 => x"ffffff",
   2384 => x"ffffff",
   2385 => x"ffffff",
   2386 => x"ffffff",
   2387 => x"ffffff",
   2388 => x"ffffff",
   2389 => x"ffffff",
   2390 => x"ffffff",
   2391 => x"ffffff",
   2392 => x"ffffff",
   2393 => x"ffffff",
   2394 => x"ffffff",
   2395 => x"ffffff",
   2396 => x"ffffff",
   2397 => x"ffffff",
   2398 => x"ffffff",
   2399 => x"ffffff",
   2400 => x"ffffff",
   2401 => x"fff540",
   2402 => x"000abf",
   2403 => x"ffffff",
   2404 => x"ffffff",
   2405 => x"fd5000",
   2406 => x"015fff",
   2407 => x"ffffff",
   2408 => x"ffffff",
   2409 => x"ffffff",
   2410 => x"ffffff",
   2411 => x"ffffff",
   2412 => x"ffffff",
   2413 => x"ffffff",
   2414 => x"ffffff",
   2415 => x"ffffff",
   2416 => x"fffffa",
   2417 => x"eb5d75",
   2418 => x"c30c30",
   2419 => x"c30c30",
   2420 => x"c30c30",
   2421 => x"c30c30",
   2422 => x"c30c30",
   2423 => x"c30c30",
   2424 => x"c30c30",
   2425 => x"c30c30",
   2426 => x"c30c30",
   2427 => x"c30c30",
   2428 => x"c30c30",
   2429 => x"d75eba",
   2430 => x"ebffff",
   2431 => x"ffffff",
   2432 => x"ffffff",
   2433 => x"ffffff",
   2434 => x"ffffff",
   2435 => x"ffffff",
   2436 => x"ffffff",
   2437 => x"ffffff",
   2438 => x"fffbae",
   2439 => x"b9d74c",
   2440 => x"30c30c",
   2441 => x"30c30c",
   2442 => x"30c30c",
   2443 => x"30c30c",
   2444 => x"30c30c",
   2445 => x"30c30c",
   2446 => x"30c30c",
   2447 => x"30c30c",
   2448 => x"30c30c",
   2449 => x"30c30c",
   2450 => x"30c31d",
   2451 => x"76ebae",
   2452 => x"ffffff",
   2453 => x"ffffff",
   2454 => x"ffffff",
   2455 => x"ffffff",
   2456 => x"ffffff",
   2457 => x"ffffff",
   2458 => x"ffffff",
   2459 => x"ffffff",
   2460 => x"ffffff",
   2461 => x"fea000",
   2462 => x"015abf",
   2463 => x"ffffff",
   2464 => x"ffffff",
   2465 => x"ffffff",
   2466 => x"ffffff",
   2467 => x"ffffff",
   2468 => x"ffffff",
   2469 => x"ffffff",
   2470 => x"ffffff",
   2471 => x"ffffff",
   2472 => x"ffffff",
   2473 => x"ffffff",
   2474 => x"ffffff",
   2475 => x"ffffff",
   2476 => x"ffffff",
   2477 => x"ffffff",
   2478 => x"ffffff",
   2479 => x"ffffff",
   2480 => x"ffffff",
   2481 => x"ffffff",
   2482 => x"ffffff",
   2483 => x"ffffff",
   2484 => x"ffffff",
   2485 => x"ffffff",
   2486 => x"ffffff",
   2487 => x"ffffff",
   2488 => x"ffffff",
   2489 => x"ffffff",
   2490 => x"ffffff",
   2491 => x"ffffff",
   2492 => x"ffffff",
   2493 => x"ffffff",
   2494 => x"ffffff",
   2495 => x"ffffff",
   2496 => x"ffffff",
   2497 => x"ffffff",
   2498 => x"ffffff",
   2499 => x"ffffff",
   2500 => x"ffffff",
   2501 => x"ffffff",
   2502 => x"ffffff",
   2503 => x"ffffff",
   2504 => x"ffffff",
   2505 => x"ffffff",
   2506 => x"ffffff",
   2507 => x"ffffea",
   2508 => x"56afff",
   2509 => x"ffffff",
   2510 => x"ffffff",
   2511 => x"ffffff",
   2512 => x"ffffff",
   2513 => x"ffffff",
   2514 => x"ffffff",
   2515 => x"ffffff",
   2516 => x"ffffff",
   2517 => x"ffffff",
   2518 => x"ffffff",
   2519 => x"ffffff",
   2520 => x"ffffff",
   2521 => x"ffffff",
   2522 => x"ffffff",
   2523 => x"ffffff",
   2524 => x"ffffff",
   2525 => x"ffffff",
   2526 => x"ffffff",
   2527 => x"ffffff",
   2528 => x"ffffff",
   2529 => x"ffffff",
   2530 => x"ffffff",
   2531 => x"ffffff",
   2532 => x"ffffff",
   2533 => x"ffffff",
   2534 => x"ffffff",
   2535 => x"ffffff",
   2536 => x"ffffff",
   2537 => x"ffffff",
   2538 => x"ffffff",
   2539 => x"ffffff",
   2540 => x"ffffff",
   2541 => x"ffffff",
   2542 => x"ffffff",
   2543 => x"ffffff",
   2544 => x"ffffff",
   2545 => x"ffffff",
   2546 => x"ffffff",
   2547 => x"ffffff",
   2548 => x"ffffff",
   2549 => x"ffffff",
   2550 => x"ffffff",
   2551 => x"ffffff",
   2552 => x"ffffff",
   2553 => x"ffffff",
   2554 => x"ffffff",
   2555 => x"ffffff",
   2556 => x"ffffff",
   2557 => x"ffffff",
   2558 => x"ffffff",
   2559 => x"ffffff",
   2560 => x"ffffff",
   2561 => x"fff540",
   2562 => x"000abf",
   2563 => x"ffffff",
   2564 => x"ffffff",
   2565 => x"fd5000",
   2566 => x"02afff",
   2567 => x"ffffff",
   2568 => x"ffffff",
   2569 => x"ffffff",
   2570 => x"ffffff",
   2571 => x"ffffff",
   2572 => x"ffffff",
   2573 => x"ffffff",
   2574 => x"ffffff",
   2575 => x"ffffff",
   2576 => x"ebad75",
   2577 => x"c30c30",
   2578 => x"c30c30",
   2579 => x"c30c30",
   2580 => x"c30c30",
   2581 => x"c30c30",
   2582 => x"c30c30",
   2583 => x"c30c30",
   2584 => x"c30c30",
   2585 => x"c30c30",
   2586 => x"c30c30",
   2587 => x"c30c30",
   2588 => x"c30c30",
   2589 => x"c30c30",
   2590 => x"d75eba",
   2591 => x"ffffff",
   2592 => x"ffffff",
   2593 => x"ffffff",
   2594 => x"ffffff",
   2595 => x"ffffff",
   2596 => x"ffffff",
   2597 => x"ffffee",
   2598 => x"b9d74c",
   2599 => x"30c30c",
   2600 => x"30c30c",
   2601 => x"30c30c",
   2602 => x"30c30c",
   2603 => x"30c30c",
   2604 => x"30c30c",
   2605 => x"30c30c",
   2606 => x"30c30c",
   2607 => x"30c30c",
   2608 => x"30c30c",
   2609 => x"30c30c",
   2610 => x"30c30c",
   2611 => x"30c31d",
   2612 => x"76ebbf",
   2613 => x"ffffff",
   2614 => x"ffffff",
   2615 => x"ffffff",
   2616 => x"ffffff",
   2617 => x"ffffff",
   2618 => x"ffffff",
   2619 => x"ffffff",
   2620 => x"ffffff",
   2621 => x"fd5000",
   2622 => x"015abf",
   2623 => x"ffffff",
   2624 => x"ffffff",
   2625 => x"ffffff",
   2626 => x"ffffff",
   2627 => x"ffffff",
   2628 => x"ffffff",
   2629 => x"ffffff",
   2630 => x"ffffff",
   2631 => x"ffffff",
   2632 => x"ffffff",
   2633 => x"ffffff",
   2634 => x"ffffff",
   2635 => x"ffffff",
   2636 => x"ffffff",
   2637 => x"ffffff",
   2638 => x"ffffff",
   2639 => x"ffffff",
   2640 => x"ffffff",
   2641 => x"ffffff",
   2642 => x"ffffff",
   2643 => x"ffffff",
   2644 => x"ffffff",
   2645 => x"ffffff",
   2646 => x"ffffff",
   2647 => x"ffffff",
   2648 => x"ffffff",
   2649 => x"ffffff",
   2650 => x"ffffff",
   2651 => x"ffffff",
   2652 => x"ffffff",
   2653 => x"ffffff",
   2654 => x"ffffff",
   2655 => x"ffffff",
   2656 => x"ffffff",
   2657 => x"ffffff",
   2658 => x"ffffff",
   2659 => x"ffffff",
   2660 => x"ffffff",
   2661 => x"ffffff",
   2662 => x"ffffff",
   2663 => x"ffffff",
   2664 => x"ffffff",
   2665 => x"ffffff",
   2666 => x"ffffff",
   2667 => x"fffa95",
   2668 => x"abffff",
   2669 => x"ffffff",
   2670 => x"ffffff",
   2671 => x"ffffff",
   2672 => x"ffffff",
   2673 => x"ffffff",
   2674 => x"ffffff",
   2675 => x"ffffff",
   2676 => x"ffffff",
   2677 => x"ffffff",
   2678 => x"ffffff",
   2679 => x"ffffff",
   2680 => x"ffffff",
   2681 => x"ffffff",
   2682 => x"ffffff",
   2683 => x"ffffff",
   2684 => x"ffffff",
   2685 => x"ffffff",
   2686 => x"ffffff",
   2687 => x"ffffff",
   2688 => x"ffffff",
   2689 => x"ffffff",
   2690 => x"ffffff",
   2691 => x"ffffff",
   2692 => x"ffffff",
   2693 => x"ffffff",
   2694 => x"ffffff",
   2695 => x"ffffff",
   2696 => x"ffffff",
   2697 => x"ffffff",
   2698 => x"ffffff",
   2699 => x"ffffff",
   2700 => x"ffffff",
   2701 => x"ffffff",
   2702 => x"ffffff",
   2703 => x"ffffff",
   2704 => x"ffffff",
   2705 => x"ffffff",
   2706 => x"ffffff",
   2707 => x"ffffff",
   2708 => x"ffffff",
   2709 => x"ffffff",
   2710 => x"ffffff",
   2711 => x"ffffff",
   2712 => x"ffffff",
   2713 => x"ffffff",
   2714 => x"ffffff",
   2715 => x"ffffff",
   2716 => x"ffffff",
   2717 => x"ffffff",
   2718 => x"ffffff",
   2719 => x"ffffff",
   2720 => x"ffffff",
   2721 => x"fff540",
   2722 => x"000abf",
   2723 => x"ffffff",
   2724 => x"ffffff",
   2725 => x"a80000",
   2726 => x"02afff",
   2727 => x"ffffff",
   2728 => x"ffffff",
   2729 => x"ffffff",
   2730 => x"ffffff",
   2731 => x"ffffff",
   2732 => x"ffffff",
   2733 => x"ffffff",
   2734 => x"ffffff",
   2735 => x"ffaeb5",
   2736 => x"c30c30",
   2737 => x"c30c30",
   2738 => x"c30c30",
   2739 => x"c30c30",
   2740 => x"c30c30",
   2741 => x"c30c30",
   2742 => x"c30c30",
   2743 => x"c30c30",
   2744 => x"c30c30",
   2745 => x"c30c30",
   2746 => x"c30c30",
   2747 => x"c30c30",
   2748 => x"c30c30",
   2749 => x"c30c30",
   2750 => x"c30c35",
   2751 => x"ebafff",
   2752 => x"ffffff",
   2753 => x"ffffff",
   2754 => x"ffffff",
   2755 => x"ffffff",
   2756 => x"ffffff",
   2757 => x"bae75d",
   2758 => x"30c30c",
   2759 => x"30c30c",
   2760 => x"30c30c",
   2761 => x"30c30c",
   2762 => x"30c30c",
   2763 => x"30c30c",
   2764 => x"30c30c",
   2765 => x"30c30c",
   2766 => x"30c30c",
   2767 => x"30c30c",
   2768 => x"30c30c",
   2769 => x"30c30c",
   2770 => x"30c30c",
   2771 => x"30c30c",
   2772 => x"30c75d",
   2773 => x"baefff",
   2774 => x"ffffff",
   2775 => x"ffffff",
   2776 => x"ffffff",
   2777 => x"ffffff",
   2778 => x"ffffff",
   2779 => x"ffffff",
   2780 => x"ffffff",
   2781 => x"fd5000",
   2782 => x"015fff",
   2783 => x"ffffff",
   2784 => x"ffffff",
   2785 => x"ffffff",
   2786 => x"ffffff",
   2787 => x"ffffff",
   2788 => x"ffffff",
   2789 => x"ffffff",
   2790 => x"ffffff",
   2791 => x"ffffff",
   2792 => x"ffffff",
   2793 => x"ffffff",
   2794 => x"ffffff",
   2795 => x"ffffff",
   2796 => x"ffffff",
   2797 => x"ffffff",
   2798 => x"ffffff",
   2799 => x"ffffff",
   2800 => x"ffffff",
   2801 => x"ffffff",
   2802 => x"ffffff",
   2803 => x"ffffff",
   2804 => x"ffffff",
   2805 => x"ffffff",
   2806 => x"ffffff",
   2807 => x"ffffff",
   2808 => x"ffffff",
   2809 => x"ffffff",
   2810 => x"ffffff",
   2811 => x"ffffff",
   2812 => x"ffffff",
   2813 => x"ffffff",
   2814 => x"ffffff",
   2815 => x"ffffff",
   2816 => x"ffffff",
   2817 => x"ffffff",
   2818 => x"ffffff",
   2819 => x"ffffff",
   2820 => x"ffffff",
   2821 => x"ffffff",
   2822 => x"ffffff",
   2823 => x"ffffff",
   2824 => x"ffffff",
   2825 => x"ffffff",
   2826 => x"ffffff",
   2827 => x"fea56a",
   2828 => x"ffffff",
   2829 => x"ffffff",
   2830 => x"ffffff",
   2831 => x"ffffff",
   2832 => x"ffffff",
   2833 => x"ffffff",
   2834 => x"ffffff",
   2835 => x"ffffff",
   2836 => x"ffffff",
   2837 => x"ffffff",
   2838 => x"ffffff",
   2839 => x"ffffff",
   2840 => x"ffffff",
   2841 => x"ffffff",
   2842 => x"ffffff",
   2843 => x"ffffff",
   2844 => x"ffffff",
   2845 => x"ffffff",
   2846 => x"ffffff",
   2847 => x"ffffff",
   2848 => x"ffffff",
   2849 => x"ffffff",
   2850 => x"ffffff",
   2851 => x"ffffff",
   2852 => x"ffffff",
   2853 => x"ffffff",
   2854 => x"ffffff",
   2855 => x"ffffff",
   2856 => x"ffffff",
   2857 => x"ffffff",
   2858 => x"ffffff",
   2859 => x"ffffff",
   2860 => x"ffffff",
   2861 => x"ffffff",
   2862 => x"ffffff",
   2863 => x"ffffff",
   2864 => x"ffffff",
   2865 => x"ffffff",
   2866 => x"ffffff",
   2867 => x"ffffff",
   2868 => x"ffffff",
   2869 => x"ffffff",
   2870 => x"ffffff",
   2871 => x"ffffff",
   2872 => x"ffffff",
   2873 => x"ffffff",
   2874 => x"ffffff",
   2875 => x"ffffff",
   2876 => x"ffffff",
   2877 => x"ffffff",
   2878 => x"ffffff",
   2879 => x"ffffff",
   2880 => x"ffffff",
   2881 => x"fff540",
   2882 => x"000abf",
   2883 => x"ffffff",
   2884 => x"ffffea",
   2885 => x"540000",
   2886 => x"57ffff",
   2887 => x"ffffff",
   2888 => x"ffffff",
   2889 => x"ffffff",
   2890 => x"ffffff",
   2891 => x"ffffff",
   2892 => x"ffffff",
   2893 => x"ffffff",
   2894 => x"fffeba",
   2895 => x"d75c30",
   2896 => x"c30c30",
   2897 => x"c30c30",
   2898 => x"c30c30",
   2899 => x"c30c30",
   2900 => x"c30c30",
   2901 => x"c30c30",
   2902 => x"c30c30",
   2903 => x"c30c30",
   2904 => x"c30c30",
   2905 => x"c30c30",
   2906 => x"c30c30",
   2907 => x"c30c30",
   2908 => x"c30c30",
   2909 => x"c30c30",
   2910 => x"c30c30",
   2911 => x"c30d7a",
   2912 => x"ebffff",
   2913 => x"ffffff",
   2914 => x"ffffff",
   2915 => x"ffffff",
   2916 => x"fffbae",
   2917 => x"74c30c",
   2918 => x"30c30c",
   2919 => x"30c30c",
   2920 => x"30c30c",
   2921 => x"30c30c",
   2922 => x"30c30c",
   2923 => x"30c30c",
   2924 => x"30c30c",
   2925 => x"30c30c",
   2926 => x"30c30c",
   2927 => x"30c30c",
   2928 => x"30c30c",
   2929 => x"30c30c",
   2930 => x"30c30c",
   2931 => x"30c30c",
   2932 => x"30c30c",
   2933 => x"31dbae",
   2934 => x"ffffff",
   2935 => x"ffffff",
   2936 => x"ffffff",
   2937 => x"ffffff",
   2938 => x"ffffff",
   2939 => x"ffffff",
   2940 => x"ffffff",
   2941 => x"fd5000",
   2942 => x"015fff",
   2943 => x"ffffff",
   2944 => x"ffffff",
   2945 => x"feaaaa",
   2946 => x"aaaaaa",
   2947 => x"aaaabf",
   2948 => x"ffffff",
   2949 => x"ffffff",
   2950 => x"ffffff",
   2951 => x"ffffff",
   2952 => x"ffffff",
   2953 => x"ffffff",
   2954 => x"ffffff",
   2955 => x"ffffff",
   2956 => x"ffffff",
   2957 => x"ffffff",
   2958 => x"ffffff",
   2959 => x"ffffff",
   2960 => x"ffffff",
   2961 => x"ffffff",
   2962 => x"ffffff",
   2963 => x"ffffff",
   2964 => x"ffffff",
   2965 => x"ffffff",
   2966 => x"ffffff",
   2967 => x"ffffff",
   2968 => x"ffffff",
   2969 => x"ffffff",
   2970 => x"ffffff",
   2971 => x"ffffff",
   2972 => x"ffffff",
   2973 => x"ffffff",
   2974 => x"ffffff",
   2975 => x"ffffff",
   2976 => x"ffffff",
   2977 => x"ffffff",
   2978 => x"ffffff",
   2979 => x"ffffff",
   2980 => x"ffffff",
   2981 => x"ffffff",
   2982 => x"ffffff",
   2983 => x"ffffff",
   2984 => x"ffffff",
   2985 => x"ffffff",
   2986 => x"ffffff",
   2987 => x"a95abf",
   2988 => x"ffffff",
   2989 => x"ffffff",
   2990 => x"ffffff",
   2991 => x"ffffff",
   2992 => x"ffffff",
   2993 => x"ffffff",
   2994 => x"ffffff",
   2995 => x"ffffff",
   2996 => x"ffffff",
   2997 => x"ffffff",
   2998 => x"ffffff",
   2999 => x"ffffff",
   3000 => x"ffffff",
   3001 => x"ffffff",
   3002 => x"ffffff",
   3003 => x"ffffff",
   3004 => x"ffffff",
   3005 => x"ffffff",
   3006 => x"ffffff",
   3007 => x"ffffff",
   3008 => x"ffffff",
   3009 => x"ffffff",
   3010 => x"ffffff",
   3011 => x"ffffff",
   3012 => x"ffffff",
   3013 => x"ffffff",
   3014 => x"ffffff",
   3015 => x"ffffff",
   3016 => x"ffffff",
   3017 => x"ffffff",
   3018 => x"ffffff",
   3019 => x"ffffff",
   3020 => x"ffffff",
   3021 => x"ffffff",
   3022 => x"ffffff",
   3023 => x"ffffff",
   3024 => x"ffffff",
   3025 => x"ffffff",
   3026 => x"ffffff",
   3027 => x"ffffff",
   3028 => x"ffffff",
   3029 => x"ffffff",
   3030 => x"ffffff",
   3031 => x"ffffff",
   3032 => x"ffffff",
   3033 => x"ffffff",
   3034 => x"ffffff",
   3035 => x"ffffff",
   3036 => x"ffffff",
   3037 => x"ffffff",
   3038 => x"ffffff",
   3039 => x"ffffff",
   3040 => x"ffffff",
   3041 => x"fff540",
   3042 => x"000abf",
   3043 => x"ffffff",
   3044 => x"fffa95",
   3045 => x"000000",
   3046 => x"abffff",
   3047 => x"ffffff",
   3048 => x"ffffff",
   3049 => x"ffffff",
   3050 => x"ffffff",
   3051 => x"ffffff",
   3052 => x"ffffff",
   3053 => x"ffffff",
   3054 => x"ebad70",
   3055 => x"c30c30",
   3056 => x"c30c30",
   3057 => x"c30c30",
   3058 => x"c30c30",
   3059 => x"c30c30",
   3060 => x"c30c30",
   3061 => x"c30c30",
   3062 => x"c30c30",
   3063 => x"c30c30",
   3064 => x"c30c30",
   3065 => x"c30c30",
   3066 => x"c30c30",
   3067 => x"c30c30",
   3068 => x"c30c30",
   3069 => x"c30c30",
   3070 => x"c30c30",
   3071 => x"c30c30",
   3072 => x"c35ebf",
   3073 => x"ffffff",
   3074 => x"ffffff",
   3075 => x"ffffee",
   3076 => x"b9d30c",
   3077 => x"30c30c",
   3078 => x"30c30c",
   3079 => x"30c30c",
   3080 => x"30c30c",
   3081 => x"30c30c",
   3082 => x"30c30c",
   3083 => x"30c30c",
   3084 => x"30c30c",
   3085 => x"30c30c",
   3086 => x"30c30c",
   3087 => x"30c30c",
   3088 => x"30c30c",
   3089 => x"30c30c",
   3090 => x"30c30c",
   3091 => x"30c30c",
   3092 => x"30c30c",
   3093 => x"30c30c",
   3094 => x"76efff",
   3095 => x"ffffff",
   3096 => x"ffffff",
   3097 => x"ffffff",
   3098 => x"ffffff",
   3099 => x"ffffff",
   3100 => x"ffffff",
   3101 => x"fd5000",
   3102 => x"015fff",
   3103 => x"ffffff",
   3104 => x"ffffff",
   3105 => x"fd5015",
   3106 => x"555555",
   3107 => x"555555",
   3108 => x"ffffff",
   3109 => x"ffffff",
   3110 => x"ffffff",
   3111 => x"ffffff",
   3112 => x"ffffff",
   3113 => x"ffffff",
   3114 => x"ffffff",
   3115 => x"ffffff",
   3116 => x"ffffff",
   3117 => x"ffffff",
   3118 => x"ffffff",
   3119 => x"ffffff",
   3120 => x"ffffff",
   3121 => x"ffffff",
   3122 => x"ffffff",
   3123 => x"ffffff",
   3124 => x"ffffff",
   3125 => x"ffffff",
   3126 => x"ffffff",
   3127 => x"ffffff",
   3128 => x"ffffff",
   3129 => x"ffffff",
   3130 => x"ffffff",
   3131 => x"ffffff",
   3132 => x"ffffff",
   3133 => x"ffffff",
   3134 => x"ffffff",
   3135 => x"ffffff",
   3136 => x"ffffff",
   3137 => x"ffffff",
   3138 => x"ffffff",
   3139 => x"ffffff",
   3140 => x"ffffff",
   3141 => x"ffffff",
   3142 => x"ffffff",
   3143 => x"ffffff",
   3144 => x"ffffff",
   3145 => x"ffffff",
   3146 => x"ffffea",
   3147 => x"56afff",
   3148 => x"ffffff",
   3149 => x"ffffff",
   3150 => x"ffffff",
   3151 => x"ffffff",
   3152 => x"ffffff",
   3153 => x"ffffff",
   3154 => x"ffffff",
   3155 => x"ffffff",
   3156 => x"ffffff",
   3157 => x"ffffff",
   3158 => x"ffffff",
   3159 => x"ffffff",
   3160 => x"ffffff",
   3161 => x"ffffff",
   3162 => x"ffffff",
   3163 => x"ffffff",
   3164 => x"ffffff",
   3165 => x"ffffff",
   3166 => x"ffffff",
   3167 => x"ffffff",
   3168 => x"ffffff",
   3169 => x"ffffff",
   3170 => x"ffffff",
   3171 => x"ffffff",
   3172 => x"ffffff",
   3173 => x"ffffff",
   3174 => x"ffffff",
   3175 => x"ffffff",
   3176 => x"ffffff",
   3177 => x"ffffff",
   3178 => x"ffffff",
   3179 => x"ffffff",
   3180 => x"ffffff",
   3181 => x"ffffff",
   3182 => x"ffffff",
   3183 => x"ffffff",
   3184 => x"ffffff",
   3185 => x"ffffff",
   3186 => x"ffffff",
   3187 => x"ffffff",
   3188 => x"ffffff",
   3189 => x"ffffff",
   3190 => x"ffffff",
   3191 => x"ffffff",
   3192 => x"ffffff",
   3193 => x"ffffff",
   3194 => x"ffffff",
   3195 => x"ffffff",
   3196 => x"ffffff",
   3197 => x"ffffff",
   3198 => x"ffffff",
   3199 => x"ffffff",
   3200 => x"ffffff",
   3201 => x"fff540",
   3202 => x"00056a",
   3203 => x"aaaaaa",
   3204 => x"555000",
   3205 => x"000015",
   3206 => x"ffffff",
   3207 => x"ffffff",
   3208 => x"ffffff",
   3209 => x"ffffff",
   3210 => x"ffffff",
   3211 => x"ffffff",
   3212 => x"ffffff",
   3213 => x"fffeba",
   3214 => x"c30c30",
   3215 => x"c30c30",
   3216 => x"c30c30",
   3217 => x"c30c30",
   3218 => x"c30c30",
   3219 => x"c30c30",
   3220 => x"c30c30",
   3221 => x"c30c30",
   3222 => x"c30c30",
   3223 => x"c30c30",
   3224 => x"c30c30",
   3225 => x"c30c30",
   3226 => x"c30c30",
   3227 => x"c30c30",
   3228 => x"c30c30",
   3229 => x"c30c30",
   3230 => x"c30c30",
   3231 => x"c30c30",
   3232 => x"c30c35",
   3233 => x"ebffff",
   3234 => x"ffffff",
   3235 => x"feeb9d",
   3236 => x"30c30c",
   3237 => x"30c30c",
   3238 => x"30c30c",
   3239 => x"30c30c",
   3240 => x"30c30c",
   3241 => x"30c30c",
   3242 => x"30c30c",
   3243 => x"30c30c",
   3244 => x"30c30c",
   3245 => x"30c30c",
   3246 => x"30c30c",
   3247 => x"30c30c",
   3248 => x"30c30c",
   3249 => x"30c30c",
   3250 => x"30c30c",
   3251 => x"30c30c",
   3252 => x"30c30c",
   3253 => x"30c30c",
   3254 => x"30c76e",
   3255 => x"ffffff",
   3256 => x"ffffff",
   3257 => x"ffffff",
   3258 => x"ffffff",
   3259 => x"ffffff",
   3260 => x"ffffff",
   3261 => x"fd5000",
   3262 => x"015fff",
   3263 => x"ffffff",
   3264 => x"ffffff",
   3265 => x"a95000",
   3266 => x"000000",
   3267 => x"000015",
   3268 => x"ffffff",
   3269 => x"ffffff",
   3270 => x"ffffff",
   3271 => x"ffffff",
   3272 => x"ffffff",
   3273 => x"ffffff",
   3274 => x"ffffff",
   3275 => x"ffffff",
   3276 => x"ffffff",
   3277 => x"ffffff",
   3278 => x"ffffff",
   3279 => x"ffffff",
   3280 => x"ffffff",
   3281 => x"ffffff",
   3282 => x"ffffff",
   3283 => x"ffffff",
   3284 => x"ffffff",
   3285 => x"ffffff",
   3286 => x"ffffff",
   3287 => x"ffffff",
   3288 => x"ffffff",
   3289 => x"ffffff",
   3290 => x"ffffff",
   3291 => x"ffffff",
   3292 => x"ffffff",
   3293 => x"ffffff",
   3294 => x"ffffff",
   3295 => x"ffffff",
   3296 => x"ffffff",
   3297 => x"ffffff",
   3298 => x"ffffff",
   3299 => x"ffffff",
   3300 => x"ffffff",
   3301 => x"ffffff",
   3302 => x"ffffff",
   3303 => x"ffffff",
   3304 => x"ffffff",
   3305 => x"ffffff",
   3306 => x"fffa95",
   3307 => x"abffff",
   3308 => x"ffffff",
   3309 => x"ffffff",
   3310 => x"ffffff",
   3311 => x"ffffff",
   3312 => x"ffffff",
   3313 => x"ffffff",
   3314 => x"ffffff",
   3315 => x"ffffff",
   3316 => x"ffffff",
   3317 => x"ffffff",
   3318 => x"ffffff",
   3319 => x"ffffff",
   3320 => x"ffffff",
   3321 => x"ffffff",
   3322 => x"ffffff",
   3323 => x"ffffff",
   3324 => x"ffffff",
   3325 => x"ffffff",
   3326 => x"ffffff",
   3327 => x"ffffff",
   3328 => x"ffffff",
   3329 => x"ffffff",
   3330 => x"ffffff",
   3331 => x"ffffff",
   3332 => x"ffffff",
   3333 => x"ffffff",
   3334 => x"ffffff",
   3335 => x"ffffff",
   3336 => x"ffffff",
   3337 => x"ffffff",
   3338 => x"ffffff",
   3339 => x"ffffff",
   3340 => x"ffffff",
   3341 => x"ffffff",
   3342 => x"ffffff",
   3343 => x"ffffff",
   3344 => x"ffffff",
   3345 => x"ffffff",
   3346 => x"ffffff",
   3347 => x"ffffff",
   3348 => x"ffffff",
   3349 => x"ffffff",
   3350 => x"ffffff",
   3351 => x"ffffff",
   3352 => x"ffffff",
   3353 => x"ffffff",
   3354 => x"ffffff",
   3355 => x"ffffff",
   3356 => x"ffffff",
   3357 => x"ffffff",
   3358 => x"ffffff",
   3359 => x"ffffff",
   3360 => x"ffffff",
   3361 => x"fff540",
   3362 => x"000000",
   3363 => x"000000",
   3364 => x"000000",
   3365 => x"01557f",
   3366 => x"ffffff",
   3367 => x"ffffff",
   3368 => x"ffffff",
   3369 => x"ffffff",
   3370 => x"ffffff",
   3371 => x"ffffff",
   3372 => x"ffffff",
   3373 => x"eb5c30",
   3374 => x"c30c30",
   3375 => x"c30c30",
   3376 => x"c30c30",
   3377 => x"c30c30",
   3378 => x"c30c30",
   3379 => x"c30c30",
   3380 => x"c30c30",
   3381 => x"c30c30",
   3382 => x"c30c30",
   3383 => x"c30c30",
   3384 => x"c30c30",
   3385 => x"c30c30",
   3386 => x"c30c30",
   3387 => x"c30c30",
   3388 => x"c30c30",
   3389 => x"c30c30",
   3390 => x"c30c30",
   3391 => x"c30c30",
   3392 => x"c30c30",
   3393 => x"c35ebf",
   3394 => x"ffffee",
   3395 => x"b9d30c",
   3396 => x"30c30c",
   3397 => x"30c30c",
   3398 => x"30c30c",
   3399 => x"30c30c",
   3400 => x"30c30c",
   3401 => x"30c30c",
   3402 => x"30c30c",
   3403 => x"30c30c",
   3404 => x"30c30c",
   3405 => x"30c30c",
   3406 => x"30c30c",
   3407 => x"30c30c",
   3408 => x"30c30c",
   3409 => x"30c30c",
   3410 => x"30c30c",
   3411 => x"30c30c",
   3412 => x"30c30c",
   3413 => x"30c30c",
   3414 => x"30c30c",
   3415 => x"76efff",
   3416 => x"ffffff",
   3417 => x"ffffff",
   3418 => x"ffffff",
   3419 => x"ffffff",
   3420 => x"ffffff",
   3421 => x"fd5000",
   3422 => x"015fff",
   3423 => x"ffffff",
   3424 => x"ffffff",
   3425 => x"fd5000",
   3426 => x"000000",
   3427 => x"000015",
   3428 => x"ffffff",
   3429 => x"ffffff",
   3430 => x"ffffff",
   3431 => x"ffffff",
   3432 => x"ffffff",
   3433 => x"ffffff",
   3434 => x"ffffff",
   3435 => x"ffffff",
   3436 => x"ffffff",
   3437 => x"ffffff",
   3438 => x"ffffff",
   3439 => x"ffffff",
   3440 => x"ffffff",
   3441 => x"ffffff",
   3442 => x"ffffff",
   3443 => x"ffffff",
   3444 => x"ffffff",
   3445 => x"ffffff",
   3446 => x"ffffff",
   3447 => x"ffffff",
   3448 => x"ffffff",
   3449 => x"ffffff",
   3450 => x"ffffff",
   3451 => x"ffffff",
   3452 => x"ffffff",
   3453 => x"ffffff",
   3454 => x"ffffff",
   3455 => x"ffffff",
   3456 => x"ffffff",
   3457 => x"ffffff",
   3458 => x"ffffff",
   3459 => x"ffffff",
   3460 => x"ffffff",
   3461 => x"ffffff",
   3462 => x"ffffff",
   3463 => x"ffffff",
   3464 => x"ffffff",
   3465 => x"ffffff",
   3466 => x"fea56a",
   3467 => x"ffffff",
   3468 => x"ffffff",
   3469 => x"ffffff",
   3470 => x"ffffff",
   3471 => x"ffffff",
   3472 => x"ffffff",
   3473 => x"ffffff",
   3474 => x"ffffff",
   3475 => x"ffffff",
   3476 => x"ffffff",
   3477 => x"ffffff",
   3478 => x"ffffff",
   3479 => x"ffffff",
   3480 => x"ffffff",
   3481 => x"ffffff",
   3482 => x"ffffff",
   3483 => x"ffffff",
   3484 => x"ffffff",
   3485 => x"ffffff",
   3486 => x"ffffff",
   3487 => x"ffffff",
   3488 => x"ffffff",
   3489 => x"ffffff",
   3490 => x"ffffff",
   3491 => x"ffffff",
   3492 => x"ffffff",
   3493 => x"ffffff",
   3494 => x"ffffff",
   3495 => x"ffffff",
   3496 => x"ffffff",
   3497 => x"ffffff",
   3498 => x"ffffff",
   3499 => x"ffffff",
   3500 => x"ffffff",
   3501 => x"ffffff",
   3502 => x"ffffff",
   3503 => x"ffffff",
   3504 => x"ffffff",
   3505 => x"ffffff",
   3506 => x"ffffff",
   3507 => x"ffffff",
   3508 => x"ffffff",
   3509 => x"ffffff",
   3510 => x"ffffff",
   3511 => x"ffffff",
   3512 => x"ffffff",
   3513 => x"ffffff",
   3514 => x"ffffff",
   3515 => x"ffffff",
   3516 => x"ffffff",
   3517 => x"ffffff",
   3518 => x"ffffff",
   3519 => x"ffffff",
   3520 => x"ffffff",
   3521 => x"fff540",
   3522 => x"000000",
   3523 => x"000000",
   3524 => x"000000",
   3525 => x"56afff",
   3526 => x"ffffff",
   3527 => x"ffffff",
   3528 => x"ffffff",
   3529 => x"ffffff",
   3530 => x"ffffff",
   3531 => x"ffffff",
   3532 => x"fffeb5",
   3533 => x"c30c30",
   3534 => x"c30c30",
   3535 => x"c30c30",
   3536 => x"c30c30",
   3537 => x"c30c30",
   3538 => x"c30c30",
   3539 => x"c30c30",
   3540 => x"c30c30",
   3541 => x"c30c30",
   3542 => x"c30c30",
   3543 => x"c30c30",
   3544 => x"c30c30",
   3545 => x"c30c30",
   3546 => x"c30c30",
   3547 => x"c30c30",
   3548 => x"c30c30",
   3549 => x"c30c30",
   3550 => x"c30c30",
   3551 => x"c30c30",
   3552 => x"c30c30",
   3553 => x"c30c35",
   3554 => x"eaeb8c",
   3555 => x"30c30c",
   3556 => x"30c30c",
   3557 => x"30c30c",
   3558 => x"30c30c",
   3559 => x"30c30c",
   3560 => x"30c30c",
   3561 => x"30c30c",
   3562 => x"30c30c",
   3563 => x"30c30c",
   3564 => x"30c30c",
   3565 => x"30c30c",
   3566 => x"30c30c",
   3567 => x"30c30c",
   3568 => x"30c30c",
   3569 => x"30c30c",
   3570 => x"30c30c",
   3571 => x"30c30c",
   3572 => x"30c30c",
   3573 => x"30c30c",
   3574 => x"30c30c",
   3575 => x"30c76e",
   3576 => x"ffffff",
   3577 => x"ffffff",
   3578 => x"ffffff",
   3579 => x"ffffff",
   3580 => x"ffffff",
   3581 => x"fd5000",
   3582 => x"015fff",
   3583 => x"ffffff",
   3584 => x"ffffff",
   3585 => x"feaaaa",
   3586 => x"aaaa95",
   3587 => x"000015",
   3588 => x"ffffff",
   3589 => x"ffffff",
   3590 => x"ffffff",
   3591 => x"ffffff",
   3592 => x"ffffff",
   3593 => x"ffffff",
   3594 => x"ffffff",
   3595 => x"ffffff",
   3596 => x"ffffff",
   3597 => x"ffffff",
   3598 => x"ffffff",
   3599 => x"ffffff",
   3600 => x"ffffff",
   3601 => x"ffffff",
   3602 => x"ffffff",
   3603 => x"ffffff",
   3604 => x"ffffff",
   3605 => x"ffffff",
   3606 => x"ffffff",
   3607 => x"ffffff",
   3608 => x"ffffff",
   3609 => x"ffffff",
   3610 => x"ffffff",
   3611 => x"ffffff",
   3612 => x"ffffff",
   3613 => x"ffffff",
   3614 => x"ffffff",
   3615 => x"ffffff",
   3616 => x"ffffff",
   3617 => x"ffffff",
   3618 => x"ffffff",
   3619 => x"ffffff",
   3620 => x"ffffff",
   3621 => x"ffffff",
   3622 => x"ffffff",
   3623 => x"ffffff",
   3624 => x"ffffff",
   3625 => x"ffffff",
   3626 => x"a95abf",
   3627 => x"ffffff",
   3628 => x"ffffff",
   3629 => x"ffffff",
   3630 => x"ffffff",
   3631 => x"ffffff",
   3632 => x"ffffff",
   3633 => x"ffffff",
   3634 => x"ffffff",
   3635 => x"ffffff",
   3636 => x"ffffff",
   3637 => x"ffffff",
   3638 => x"ffffff",
   3639 => x"ffffff",
   3640 => x"ffffff",
   3641 => x"ffffff",
   3642 => x"ffffff",
   3643 => x"ffffff",
   3644 => x"ffffff",
   3645 => x"ffffff",
   3646 => x"ffffff",
   3647 => x"ffffff",
   3648 => x"ffffff",
   3649 => x"ffffff",
   3650 => x"ffffff",
   3651 => x"ffffff",
   3652 => x"ffffff",
   3653 => x"ffffff",
   3654 => x"ffffff",
   3655 => x"ffffff",
   3656 => x"ffffff",
   3657 => x"ffffff",
   3658 => x"ffffff",
   3659 => x"ffffff",
   3660 => x"ffffff",
   3661 => x"ffffff",
   3662 => x"ffffff",
   3663 => x"ffffff",
   3664 => x"ffffff",
   3665 => x"ffffff",
   3666 => x"ffffff",
   3667 => x"ffffff",
   3668 => x"ffffff",
   3669 => x"ffffff",
   3670 => x"ffffff",
   3671 => x"ffffff",
   3672 => x"ffffff",
   3673 => x"ffffff",
   3674 => x"ffffff",
   3675 => x"ffffff",
   3676 => x"ffffff",
   3677 => x"ffffff",
   3678 => x"ffffff",
   3679 => x"ffffff",
   3680 => x"ffffff",
   3681 => x"fff540",
   3682 => x"000015",
   3683 => x"555540",
   3684 => x"000000",
   3685 => x"015abf",
   3686 => x"ffffff",
   3687 => x"ffffff",
   3688 => x"ffffff",
   3689 => x"ffffff",
   3690 => x"ffffff",
   3691 => x"ffffff",
   3692 => x"eb5c30",
   3693 => x"c30c30",
   3694 => x"c30c30",
   3695 => x"c30c30",
   3696 => x"c30c30",
   3697 => x"c30c30",
   3698 => x"c30c30",
   3699 => x"c30c30",
   3700 => x"c30c30",
   3701 => x"c30c30",
   3702 => x"c30c30",
   3703 => x"c30c30",
   3704 => x"c30c30",
   3705 => x"c30c30",
   3706 => x"c30c30",
   3707 => x"c30c30",
   3708 => x"c30c30",
   3709 => x"c30c30",
   3710 => x"c30c30",
   3711 => x"c30c30",
   3712 => x"c30c30",
   3713 => x"c30c30",
   3714 => x"a1c30c",
   3715 => x"30c30c",
   3716 => x"30c30c",
   3717 => x"30c30c",
   3718 => x"30c30c",
   3719 => x"30c30c",
   3720 => x"30c30c",
   3721 => x"30c30c",
   3722 => x"30c30c",
   3723 => x"30c30c",
   3724 => x"30c30c",
   3725 => x"30c30c",
   3726 => x"30c30c",
   3727 => x"30c30c",
   3728 => x"30c30c",
   3729 => x"30c30c",
   3730 => x"30c30c",
   3731 => x"30c30c",
   3732 => x"30c30c",
   3733 => x"30c30c",
   3734 => x"30c30c",
   3735 => x"30c30c",
   3736 => x"76efff",
   3737 => x"ffffff",
   3738 => x"ffffff",
   3739 => x"ffffff",
   3740 => x"ffffff",
   3741 => x"fea000",
   3742 => x"015abf",
   3743 => x"ffffff",
   3744 => x"ffffff",
   3745 => x"ffffff",
   3746 => x"ffffea",
   3747 => x"000015",
   3748 => x"ffffff",
   3749 => x"ffffff",
   3750 => x"ffffff",
   3751 => x"ffffff",
   3752 => x"ffffff",
   3753 => x"ffffff",
   3754 => x"ffffff",
   3755 => x"ffffff",
   3756 => x"ffffff",
   3757 => x"ffffff",
   3758 => x"ffffff",
   3759 => x"ffffff",
   3760 => x"ffffff",
   3761 => x"ffffff",
   3762 => x"ffffff",
   3763 => x"ffffff",
   3764 => x"ffffff",
   3765 => x"ffffff",
   3766 => x"ffffff",
   3767 => x"ffffff",
   3768 => x"ffffff",
   3769 => x"ffffff",
   3770 => x"ffffff",
   3771 => x"ffffff",
   3772 => x"ffffff",
   3773 => x"ffffff",
   3774 => x"ffffff",
   3775 => x"ffffff",
   3776 => x"ffffff",
   3777 => x"ffffff",
   3778 => x"ffffff",
   3779 => x"ffffff",
   3780 => x"ffffff",
   3781 => x"ffffff",
   3782 => x"ffffff",
   3783 => x"ffffff",
   3784 => x"ffffff",
   3785 => x"ffffea",
   3786 => x"56afff",
   3787 => x"ffffff",
   3788 => x"ffffff",
   3789 => x"ffffff",
   3790 => x"ffffff",
   3791 => x"ffffff",
   3792 => x"ffffff",
   3793 => x"ffffff",
   3794 => x"ffffff",
   3795 => x"ffffff",
   3796 => x"ffffff",
   3797 => x"ffffff",
   3798 => x"ffffff",
   3799 => x"ffffff",
   3800 => x"ffffff",
   3801 => x"ffffff",
   3802 => x"ffffff",
   3803 => x"ffffff",
   3804 => x"ffffff",
   3805 => x"ffffff",
   3806 => x"ffffff",
   3807 => x"ffffff",
   3808 => x"ffffff",
   3809 => x"ffffff",
   3810 => x"ffffff",
   3811 => x"ffffff",
   3812 => x"ffffff",
   3813 => x"ffffff",
   3814 => x"ffffff",
   3815 => x"ffffff",
   3816 => x"ffffff",
   3817 => x"ffffff",
   3818 => x"ffffff",
   3819 => x"ffffff",
   3820 => x"ffffff",
   3821 => x"ffffff",
   3822 => x"ffffff",
   3823 => x"ffffff",
   3824 => x"ffffff",
   3825 => x"ffffff",
   3826 => x"ffffff",
   3827 => x"ffffff",
   3828 => x"ffffff",
   3829 => x"ffffff",
   3830 => x"ffffff",
   3831 => x"ffffff",
   3832 => x"ffffff",
   3833 => x"ffffff",
   3834 => x"ffffff",
   3835 => x"ffffff",
   3836 => x"ffffff",
   3837 => x"ffffff",
   3838 => x"ffffff",
   3839 => x"ffffff",
   3840 => x"ffffff",
   3841 => x"fff540",
   3842 => x"000abf",
   3843 => x"ffffff",
   3844 => x"fea540",
   3845 => x"00002a",
   3846 => x"ffffff",
   3847 => x"ffffff",
   3848 => x"ffffff",
   3849 => x"ffffff",
   3850 => x"ffffff",
   3851 => x"fffffa",
   3852 => x"c30c30",
   3853 => x"c30c30",
   3854 => x"c30c30",
   3855 => x"c30c30",
   3856 => x"c30c30",
   3857 => x"c30c30",
   3858 => x"c30c30",
   3859 => x"c30c30",
   3860 => x"c30c30",
   3861 => x"c30c30",
   3862 => x"c30c30",
   3863 => x"c30c30",
   3864 => x"c30c30",
   3865 => x"c30c30",
   3866 => x"c30c30",
   3867 => x"c30c30",
   3868 => x"c30c30",
   3869 => x"c30c30",
   3870 => x"c30c30",
   3871 => x"c30c30",
   3872 => x"c30c30",
   3873 => x"c30918",
   3874 => x"b2c70c",
   3875 => x"30c30c",
   3876 => x"30c30c",
   3877 => x"30c30c",
   3878 => x"30c30c",
   3879 => x"30c30c",
   3880 => x"30c30c",
   3881 => x"30c30c",
   3882 => x"30c30c",
   3883 => x"30c30c",
   3884 => x"30c30c",
   3885 => x"30c30c",
   3886 => x"30c30c",
   3887 => x"30c30c",
   3888 => x"30c30c",
   3889 => x"30c30c",
   3890 => x"30c30c",
   3891 => x"30c30c",
   3892 => x"30c30c",
   3893 => x"30c30c",
   3894 => x"30c30c",
   3895 => x"30c30c",
   3896 => x"30c76e",
   3897 => x"ffffff",
   3898 => x"ffffff",
   3899 => x"ffffff",
   3900 => x"ffffff",
   3901 => x"fea000",
   3902 => x"000abf",
   3903 => x"ffffff",
   3904 => x"ffffff",
   3905 => x"ffffff",
   3906 => x"ffffea",
   3907 => x"000015",
   3908 => x"ffffff",
   3909 => x"ffffff",
   3910 => x"ffffff",
   3911 => x"ffffff",
   3912 => x"ffffff",
   3913 => x"ffffff",
   3914 => x"ffffff",
   3915 => x"ffffff",
   3916 => x"ffffff",
   3917 => x"ffffff",
   3918 => x"ffffff",
   3919 => x"ffffff",
   3920 => x"ffffff",
   3921 => x"ffffff",
   3922 => x"ffffff",
   3923 => x"ffffff",
   3924 => x"ffffff",
   3925 => x"ffffff",
   3926 => x"ffffff",
   3927 => x"ffffff",
   3928 => x"ffffff",
   3929 => x"ffffff",
   3930 => x"ffffff",
   3931 => x"ffffff",
   3932 => x"ffffff",
   3933 => x"ffffff",
   3934 => x"ffffff",
   3935 => x"ffffff",
   3936 => x"ffffff",
   3937 => x"ffffff",
   3938 => x"ffffff",
   3939 => x"ffffff",
   3940 => x"ffffff",
   3941 => x"ffffff",
   3942 => x"ffffff",
   3943 => x"ffffff",
   3944 => x"ffffff",
   3945 => x"fffa95",
   3946 => x"abffff",
   3947 => x"ffffff",
   3948 => x"ffffff",
   3949 => x"ffffff",
   3950 => x"ffffff",
   3951 => x"ffffff",
   3952 => x"ffffff",
   3953 => x"ffffff",
   3954 => x"ffffff",
   3955 => x"ffffff",
   3956 => x"ffffff",
   3957 => x"ffffff",
   3958 => x"ffffff",
   3959 => x"ffffff",
   3960 => x"ffffff",
   3961 => x"ffffff",
   3962 => x"ffffff",
   3963 => x"ffffff",
   3964 => x"ffffff",
   3965 => x"ffffff",
   3966 => x"ffffff",
   3967 => x"ffffff",
   3968 => x"ffffff",
   3969 => x"ffffff",
   3970 => x"ffffff",
   3971 => x"ffffff",
   3972 => x"ffffff",
   3973 => x"ffffff",
   3974 => x"ffffff",
   3975 => x"ffffff",
   3976 => x"ffffff",
   3977 => x"ffffff",
   3978 => x"ffffff",
   3979 => x"ffffff",
   3980 => x"ffffff",
   3981 => x"ffffff",
   3982 => x"ffffff",
   3983 => x"ffffff",
   3984 => x"ffffff",
   3985 => x"ffffff",
   3986 => x"ffffff",
   3987 => x"ffffff",
   3988 => x"ffffff",
   3989 => x"ffffff",
   3990 => x"ffffff",
   3991 => x"ffffff",
   3992 => x"ffffff",
   3993 => x"ffffff",
   3994 => x"ffffff",
   3995 => x"ffffff",
   3996 => x"ffffff",
   3997 => x"ffffff",
   3998 => x"ffffff",
   3999 => x"ffffff",
   4000 => x"ffffff",
   4001 => x"fff540",
   4002 => x"000abf",
   4003 => x"ffffff",
   4004 => x"fffa95",
   4005 => x"000015",
   4006 => x"ffffff",
   4007 => x"ffffff",
   4008 => x"ffffff",
   4009 => x"ffffff",
   4010 => x"ffffff",
   4011 => x"ffad70",
   4012 => x"c30c30",
   4013 => x"c30c30",
   4014 => x"c30c30",
   4015 => x"c30c30",
   4016 => x"c30c30",
   4017 => x"c30c30",
   4018 => x"c30c30",
   4019 => x"c30c30",
   4020 => x"c30c30",
   4021 => x"c30c30",
   4022 => x"c30c30",
   4023 => x"c30c30",
   4024 => x"c30c30",
   4025 => x"c30c30",
   4026 => x"c30c30",
   4027 => x"c30c30",
   4028 => x"c30c30",
   4029 => x"c30c30",
   4030 => x"c30c30",
   4031 => x"c30c30",
   4032 => x"c30c30",
   4033 => x"d28b3c",
   4034 => x"f3cf2c",
   4035 => x"70c30c",
   4036 => x"30c30c",
   4037 => x"30c30c",
   4038 => x"30c30c",
   4039 => x"30c30c",
   4040 => x"30c30c",
   4041 => x"30c30c",
   4042 => x"30c30c",
   4043 => x"30c30c",
   4044 => x"30c30c",
   4045 => x"30c30c",
   4046 => x"30c30c",
   4047 => x"30c30c",
   4048 => x"30c30c",
   4049 => x"30c30c",
   4050 => x"30c30c",
   4051 => x"30c30c",
   4052 => x"30c30c",
   4053 => x"30c30c",
   4054 => x"30c30c",
   4055 => x"30c30c",
   4056 => x"30c30c",
   4057 => x"77ffff",
   4058 => x"ffffff",
   4059 => x"ffffff",
   4060 => x"ffffff",
   4061 => x"fff540",
   4062 => x"000abf",
   4063 => x"ffffff",
   4064 => x"ffffff",
   4065 => x"ffffff",
   4066 => x"ffffea",
   4067 => x"000015",
   4068 => x"ffffff",
   4069 => x"ffffff",
   4070 => x"ffffff",
   4071 => x"ffffff",
   4072 => x"ffffff",
   4073 => x"ffffff",
   4074 => x"ffffff",
   4075 => x"ffffff",
   4076 => x"ffffff",
   4077 => x"ffffff",
   4078 => x"ffffff",
   4079 => x"ffffff",
   4080 => x"ffffff",
   4081 => x"ffffff",
   4082 => x"ffffff",
   4083 => x"ffffff",
   4084 => x"ffffff",
   4085 => x"ffffff",
   4086 => x"ffffff",
   4087 => x"ffffff",
   4088 => x"ffffff",
   4089 => x"ffffff",
   4090 => x"ffffff",
   4091 => x"ffffff",
   4092 => x"ffffff",
   4093 => x"ffffff",
   4094 => x"ffffff",
   4095 => x"ffffff",
   4096 => x"ffffff",
   4097 => x"ffffff",
   4098 => x"ffffff",
   4099 => x"ffffff",
   4100 => x"ffffff",
   4101 => x"ffffff",
   4102 => x"ffffff",
   4103 => x"ffffff",
   4104 => x"ffffff",
   4105 => x"fea56a",
   4106 => x"ffffff",
   4107 => x"ffffff",
   4108 => x"ffffff",
   4109 => x"ffffff",
   4110 => x"ffffff",
   4111 => x"ffffff",
   4112 => x"ffffff",
   4113 => x"ffffff",
   4114 => x"ffffff",
   4115 => x"ffffff",
   4116 => x"ffffff",
   4117 => x"ffffff",
   4118 => x"ffffff",
   4119 => x"ffffff",
   4120 => x"ffffff",
   4121 => x"ffffff",
   4122 => x"ffffff",
   4123 => x"ffffff",
   4124 => x"ffffff",
   4125 => x"ffffff",
   4126 => x"ffffff",
   4127 => x"ffffff",
   4128 => x"ffffff",
   4129 => x"ffffff",
   4130 => x"ffffff",
   4131 => x"ffffff",
   4132 => x"ffffff",
   4133 => x"ffffff",
   4134 => x"ffffff",
   4135 => x"ffffff",
   4136 => x"ffffff",
   4137 => x"ffffff",
   4138 => x"ffffff",
   4139 => x"ffffff",
   4140 => x"ffffff",
   4141 => x"ffffff",
   4142 => x"ffffff",
   4143 => x"ffffff",
   4144 => x"ffffff",
   4145 => x"ffffff",
   4146 => x"ffffff",
   4147 => x"ffffff",
   4148 => x"ffffff",
   4149 => x"ffffff",
   4150 => x"ffffff",
   4151 => x"ffffff",
   4152 => x"ffffff",
   4153 => x"ffffff",
   4154 => x"ffffff",
   4155 => x"ffffff",
   4156 => x"ffffff",
   4157 => x"ffffff",
   4158 => x"ffffff",
   4159 => x"ffffff",
   4160 => x"ffffff",
   4161 => x"fff540",
   4162 => x"000abf",
   4163 => x"ffffff",
   4164 => x"ffffea",
   4165 => x"540000",
   4166 => x"57ffff",
   4167 => x"ffffff",
   4168 => x"ffffff",
   4169 => x"ffffff",
   4170 => x"fffffa",
   4171 => x"d70c30",
   4172 => x"c30c30",
   4173 => x"c30c30",
   4174 => x"c30c30",
   4175 => x"c30c30",
   4176 => x"c30c30",
   4177 => x"c30c30",
   4178 => x"c30c30",
   4179 => x"c30c30",
   4180 => x"c30c30",
   4181 => x"c30c30",
   4182 => x"c30c30",
   4183 => x"c30c30",
   4184 => x"c30c30",
   4185 => x"c30c30",
   4186 => x"c30c30",
   4187 => x"c30c30",
   4188 => x"c30c30",
   4189 => x"c30c30",
   4190 => x"c30c30",
   4191 => x"c30c30",
   4192 => x"c30c24",
   4193 => x"b3cf3c",
   4194 => x"f3cf3c",
   4195 => x"f2c70c",
   4196 => x"30c30c",
   4197 => x"30c30c",
   4198 => x"30c30c",
   4199 => x"30c30c",
   4200 => x"30c30c",
   4201 => x"30c30c",
   4202 => x"30c30c",
   4203 => x"30c30c",
   4204 => x"30c30c",
   4205 => x"30c30c",
   4206 => x"30c30c",
   4207 => x"30c30c",
   4208 => x"30c30c",
   4209 => x"30c30c",
   4210 => x"30c30c",
   4211 => x"30c30c",
   4212 => x"30c30c",
   4213 => x"30c30c",
   4214 => x"30c30c",
   4215 => x"30c30c",
   4216 => x"30c30c",
   4217 => x"31dbbf",
   4218 => x"ffffff",
   4219 => x"ffffff",
   4220 => x"ffffff",
   4221 => x"fff540",
   4222 => x"00056a",
   4223 => x"ffffff",
   4224 => x"ffffff",
   4225 => x"ffffff",
   4226 => x"ffffea",
   4227 => x"000015",
   4228 => x"ffffff",
   4229 => x"ffffff",
   4230 => x"ffffff",
   4231 => x"ffffff",
   4232 => x"ffffff",
   4233 => x"ffffff",
   4234 => x"ffffff",
   4235 => x"ffffff",
   4236 => x"ffffff",
   4237 => x"ffffff",
   4238 => x"ffffff",
   4239 => x"ffffff",
   4240 => x"ffffff",
   4241 => x"ffffff",
   4242 => x"ffffff",
   4243 => x"ffffff",
   4244 => x"ffffff",
   4245 => x"ffffff",
   4246 => x"ffffff",
   4247 => x"ffffff",
   4248 => x"ffffff",
   4249 => x"ffffff",
   4250 => x"ffffff",
   4251 => x"ffffff",
   4252 => x"ffffff",
   4253 => x"ffffff",
   4254 => x"ffffff",
   4255 => x"ffffff",
   4256 => x"ffffff",
   4257 => x"ffffff",
   4258 => x"ffffff",
   4259 => x"ffffff",
   4260 => x"ffffff",
   4261 => x"ffffff",
   4262 => x"ffffff",
   4263 => x"ffffff",
   4264 => x"ffffff",
   4265 => x"a95abf",
   4266 => x"ffffff",
   4267 => x"ffffff",
   4268 => x"ffffff",
   4269 => x"ffffff",
   4270 => x"ffffff",
   4271 => x"ffffff",
   4272 => x"ffffff",
   4273 => x"ffffff",
   4274 => x"ffffff",
   4275 => x"ffffff",
   4276 => x"ffffff",
   4277 => x"ffffff",
   4278 => x"ffffff",
   4279 => x"ffffff",
   4280 => x"ffffff",
   4281 => x"ffffff",
   4282 => x"ffffff",
   4283 => x"ffffff",
   4284 => x"ffffff",
   4285 => x"ffffff",
   4286 => x"ffffff",
   4287 => x"ffffff",
   4288 => x"ffffff",
   4289 => x"ffffff",
   4290 => x"ffffff",
   4291 => x"ffffff",
   4292 => x"ffffff",
   4293 => x"ffffff",
   4294 => x"ffffff",
   4295 => x"ffffff",
   4296 => x"ffffff",
   4297 => x"ffffff",
   4298 => x"ffffff",
   4299 => x"ffffff",
   4300 => x"ffffff",
   4301 => x"ffffff",
   4302 => x"ffffff",
   4303 => x"ffffff",
   4304 => x"ffffff",
   4305 => x"ffffff",
   4306 => x"ffffff",
   4307 => x"ffffff",
   4308 => x"ffffff",
   4309 => x"ffffff",
   4310 => x"ffffff",
   4311 => x"ffffff",
   4312 => x"ffffff",
   4313 => x"ffffff",
   4314 => x"ffffff",
   4315 => x"ffffff",
   4316 => x"ffffff",
   4317 => x"ffffff",
   4318 => x"ffffff",
   4319 => x"ffffff",
   4320 => x"ffffff",
   4321 => x"fff540",
   4322 => x"000abf",
   4323 => x"ffffff",
   4324 => x"ffffff",
   4325 => x"a80000",
   4326 => x"02afff",
   4327 => x"ffffff",
   4328 => x"ffffff",
   4329 => x"ffffff",
   4330 => x"fffeb5",
   4331 => x"c30c30",
   4332 => x"c30c30",
   4333 => x"c30c30",
   4334 => x"c30c30",
   4335 => x"c30c30",
   4336 => x"c30c30",
   4337 => x"c30c30",
   4338 => x"c30c30",
   4339 => x"c30c30",
   4340 => x"c30c30",
   4341 => x"c30c30",
   4342 => x"c30c30",
   4343 => x"c30c30",
   4344 => x"c30c30",
   4345 => x"c30c30",
   4346 => x"c30c30",
   4347 => x"c30c30",
   4348 => x"c30c30",
   4349 => x"c30c30",
   4350 => x"c30c30",
   4351 => x"c30c30",
   4352 => x"c2462c",
   4353 => x"f3cf3c",
   4354 => x"f3cf3c",
   4355 => x"f3cf2c",
   4356 => x"70c30c",
   4357 => x"30c30c",
   4358 => x"30c30c",
   4359 => x"30c30c",
   4360 => x"30c30c",
   4361 => x"30c30c",
   4362 => x"30c30c",
   4363 => x"30c30c",
   4364 => x"30c30c",
   4365 => x"30c30c",
   4366 => x"30c30c",
   4367 => x"30c30c",
   4368 => x"30c30c",
   4369 => x"30c30c",
   4370 => x"30c30c",
   4371 => x"30c30c",
   4372 => x"30c30c",
   4373 => x"30c30c",
   4374 => x"30c30c",
   4375 => x"30c30c",
   4376 => x"30c30c",
   4377 => x"30c31d",
   4378 => x"bbffff",
   4379 => x"ffffff",
   4380 => x"ffffff",
   4381 => x"fffa80",
   4382 => x"00002a",
   4383 => x"ffffff",
   4384 => x"ffffff",
   4385 => x"ffffff",
   4386 => x"ffffea",
   4387 => x"000015",
   4388 => x"ffffff",
   4389 => x"ffffff",
   4390 => x"ffffff",
   4391 => x"ffffff",
   4392 => x"ffffff",
   4393 => x"ffffff",
   4394 => x"ffffff",
   4395 => x"ffffff",
   4396 => x"ffffff",
   4397 => x"ffffff",
   4398 => x"ffffff",
   4399 => x"ffffff",
   4400 => x"ffffff",
   4401 => x"ffffff",
   4402 => x"ffffff",
   4403 => x"ffffff",
   4404 => x"ffffff",
   4405 => x"ffffff",
   4406 => x"ffffff",
   4407 => x"ffffff",
   4408 => x"ffffff",
   4409 => x"ffffff",
   4410 => x"ffffff",
   4411 => x"ffffff",
   4412 => x"ffffff",
   4413 => x"ffffff",
   4414 => x"ffffff",
   4415 => x"ffffff",
   4416 => x"ffffff",
   4417 => x"ffffff",
   4418 => x"ffffff",
   4419 => x"ffffff",
   4420 => x"ffffff",
   4421 => x"ffffff",
   4422 => x"ffffff",
   4423 => x"ffffff",
   4424 => x"ffffea",
   4425 => x"56afff",
   4426 => x"ffffff",
   4427 => x"ffffff",
   4428 => x"ffffff",
   4429 => x"ffffff",
   4430 => x"ffffff",
   4431 => x"ffffff",
   4432 => x"ffffff",
   4433 => x"ffffff",
   4434 => x"ffffff",
   4435 => x"ffffff",
   4436 => x"ffffff",
   4437 => x"ffffff",
   4438 => x"ffffff",
   4439 => x"ffffff",
   4440 => x"ffffff",
   4441 => x"ffffff",
   4442 => x"ffffff",
   4443 => x"ffffff",
   4444 => x"ffffff",
   4445 => x"ffffff",
   4446 => x"ffffff",
   4447 => x"ffffff",
   4448 => x"ffffff",
   4449 => x"ffffff",
   4450 => x"ffffff",
   4451 => x"ffffff",
   4452 => x"ffffff",
   4453 => x"ffffff",
   4454 => x"ffffff",
   4455 => x"ffffff",
   4456 => x"ffffff",
   4457 => x"ffffff",
   4458 => x"ffffff",
   4459 => x"ffffff",
   4460 => x"ffffff",
   4461 => x"ffffff",
   4462 => x"ffffff",
   4463 => x"ffffff",
   4464 => x"ffffff",
   4465 => x"ffffff",
   4466 => x"ffffff",
   4467 => x"ffffff",
   4468 => x"ffffff",
   4469 => x"ffffff",
   4470 => x"ffffff",
   4471 => x"ffffff",
   4472 => x"ffffff",
   4473 => x"ffffff",
   4474 => x"ffffff",
   4475 => x"ffffff",
   4476 => x"ffffff",
   4477 => x"ffffff",
   4478 => x"ffffff",
   4479 => x"ffffff",
   4480 => x"ffffff",
   4481 => x"fff540",
   4482 => x"000abf",
   4483 => x"ffffff",
   4484 => x"ffffff",
   4485 => x"fd5000",
   4486 => x"015fff",
   4487 => x"ffffff",
   4488 => x"ffffff",
   4489 => x"ffffff",
   4490 => x"eb5c30",
   4491 => x"c30c30",
   4492 => x"c30c30",
   4493 => x"c30c30",
   4494 => x"c30c30",
   4495 => x"c30c30",
   4496 => x"c30c30",
   4497 => x"c30c30",
   4498 => x"c30c30",
   4499 => x"c30c30",
   4500 => x"c30c30",
   4501 => x"c30c30",
   4502 => x"c30c30",
   4503 => x"c30c30",
   4504 => x"c30c30",
   4505 => x"c30c30",
   4506 => x"c30c30",
   4507 => x"c30c30",
   4508 => x"c30c30",
   4509 => x"c30c30",
   4510 => x"c30c30",
   4511 => x"c30c30",
   4512 => x"a2cf3c",
   4513 => x"f3cf3c",
   4514 => x"f3cf3c",
   4515 => x"f3cf3c",
   4516 => x"b1c30c",
   4517 => x"30c30c",
   4518 => x"30c30c",
   4519 => x"30c30c",
   4520 => x"30c30c",
   4521 => x"30c30c",
   4522 => x"30c30c",
   4523 => x"30c30c",
   4524 => x"30c30c",
   4525 => x"30c30c",
   4526 => x"30c30c",
   4527 => x"30c30c",
   4528 => x"30c30c",
   4529 => x"30c30c",
   4530 => x"30c30c",
   4531 => x"30c30c",
   4532 => x"30c30c",
   4533 => x"30c30c",
   4534 => x"30c30c",
   4535 => x"30c30c",
   4536 => x"30c30c",
   4537 => x"30c30c",
   4538 => x"32efff",
   4539 => x"ffffff",
   4540 => x"ffffff",
   4541 => x"ffffd5",
   4542 => x"000015",
   4543 => x"abffff",
   4544 => x"ffffff",
   4545 => x"ffffff",
   4546 => x"ffffea",
   4547 => x"000015",
   4548 => x"ffffff",
   4549 => x"ffffff",
   4550 => x"ffffff",
   4551 => x"ffffff",
   4552 => x"ffffff",
   4553 => x"ffffff",
   4554 => x"ffffff",
   4555 => x"ffffff",
   4556 => x"ffffff",
   4557 => x"ffffff",
   4558 => x"ffffff",
   4559 => x"ffffff",
   4560 => x"ffffff",
   4561 => x"ffffff",
   4562 => x"ffffff",
   4563 => x"ffffff",
   4564 => x"ffffff",
   4565 => x"ffffff",
   4566 => x"ffffff",
   4567 => x"ffffff",
   4568 => x"ffffff",
   4569 => x"ffffff",
   4570 => x"ffffff",
   4571 => x"ffffff",
   4572 => x"ffffff",
   4573 => x"ffffff",
   4574 => x"ffffff",
   4575 => x"ffffff",
   4576 => x"ffffff",
   4577 => x"ffffff",
   4578 => x"ffffff",
   4579 => x"ffffff",
   4580 => x"ffffff",
   4581 => x"ffffff",
   4582 => x"ffffff",
   4583 => x"ffffff",
   4584 => x"fffa95",
   4585 => x"abffff",
   4586 => x"ffffff",
   4587 => x"ffffff",
   4588 => x"ffffff",
   4589 => x"ffffff",
   4590 => x"ffffff",
   4591 => x"ffffff",
   4592 => x"ffffff",
   4593 => x"ffffff",
   4594 => x"ffffff",
   4595 => x"ffffff",
   4596 => x"ffffff",
   4597 => x"ffffff",
   4598 => x"ffffff",
   4599 => x"ffffff",
   4600 => x"ffffff",
   4601 => x"ffffff",
   4602 => x"ffffff",
   4603 => x"ffffff",
   4604 => x"ffffff",
   4605 => x"ffffff",
   4606 => x"ffffff",
   4607 => x"ffffff",
   4608 => x"ffffff",
   4609 => x"ffffff",
   4610 => x"ffffff",
   4611 => x"ffffff",
   4612 => x"ffffff",
   4613 => x"ffffff",
   4614 => x"ffffff",
   4615 => x"ffffff",
   4616 => x"ffffff",
   4617 => x"ffffff",
   4618 => x"ffffff",
   4619 => x"ffffff",
   4620 => x"ffffff",
   4621 => x"ffffff",
   4622 => x"ffffff",
   4623 => x"ffffff",
   4624 => x"ffffff",
   4625 => x"ffffff",
   4626 => x"ffffff",
   4627 => x"ffffff",
   4628 => x"ffffff",
   4629 => x"ffffff",
   4630 => x"ffffff",
   4631 => x"ffffff",
   4632 => x"ffffff",
   4633 => x"ffffff",
   4634 => x"ffffff",
   4635 => x"ffffff",
   4636 => x"ffffff",
   4637 => x"ffffff",
   4638 => x"ffffff",
   4639 => x"ffffff",
   4640 => x"ffffff",
   4641 => x"fff540",
   4642 => x"000abf",
   4643 => x"ffffff",
   4644 => x"ffffff",
   4645 => x"fea000",
   4646 => x"000abf",
   4647 => x"ffffff",
   4648 => x"ffffff",
   4649 => x"fffffa",
   4650 => x"d70c30",
   4651 => x"c30c30",
   4652 => x"c30c30",
   4653 => x"c30c30",
   4654 => x"c30c30",
   4655 => x"c30c30",
   4656 => x"c30c30",
   4657 => x"c30c30",
   4658 => x"c30c30",
   4659 => x"c30c30",
   4660 => x"c30c30",
   4661 => x"c30c30",
   4662 => x"c30c30",
   4663 => x"c30c30",
   4664 => x"c30c30",
   4665 => x"c30c30",
   4666 => x"c30c30",
   4667 => x"c30c30",
   4668 => x"c30c30",
   4669 => x"c30c30",
   4670 => x"c30c30",
   4671 => x"c30918",
   4672 => x"b3cf3c",
   4673 => x"f3cf3c",
   4674 => x"f3cf3c",
   4675 => x"f3cf3c",
   4676 => x"f3cb0c",
   4677 => x"30c30c",
   4678 => x"30c30c",
   4679 => x"30c30c",
   4680 => x"30c30c",
   4681 => x"30c30c",
   4682 => x"30c30c",
   4683 => x"30c30c",
   4684 => x"30c30c",
   4685 => x"30c30c",
   4686 => x"30c30c",
   4687 => x"30c30c",
   4688 => x"30c30c",
   4689 => x"30c30c",
   4690 => x"30c30c",
   4691 => x"30c30c",
   4692 => x"30c30c",
   4693 => x"30c30c",
   4694 => x"30c30c",
   4695 => x"30c30c",
   4696 => x"30c30c",
   4697 => x"30c30c",
   4698 => x"30c77f",
   4699 => x"ffffff",
   4700 => x"ffffff",
   4701 => x"ffffea",
   4702 => x"540000",
   4703 => x"56afff",
   4704 => x"ffffff",
   4705 => x"ffffff",
   4706 => x"ffffea",
   4707 => x"000015",
   4708 => x"ffffff",
   4709 => x"ffffff",
   4710 => x"ffffff",
   4711 => x"ffffff",
   4712 => x"ffffff",
   4713 => x"ffffff",
   4714 => x"ffffff",
   4715 => x"ffffff",
   4716 => x"ffffff",
   4717 => x"ffffff",
   4718 => x"ffffff",
   4719 => x"ffffff",
   4720 => x"ffffff",
   4721 => x"ffffff",
   4722 => x"ffffff",
   4723 => x"ffffff",
   4724 => x"ffffff",
   4725 => x"ffffff",
   4726 => x"ffffff",
   4727 => x"ffffff",
   4728 => x"ffffff",
   4729 => x"ffffff",
   4730 => x"ffffff",
   4731 => x"ffffff",
   4732 => x"ffffff",
   4733 => x"ffffff",
   4734 => x"ffffff",
   4735 => x"ffffff",
   4736 => x"ffffff",
   4737 => x"ffffff",
   4738 => x"ffffff",
   4739 => x"ffffff",
   4740 => x"ffffff",
   4741 => x"ffffff",
   4742 => x"ffffff",
   4743 => x"ffffff",
   4744 => x"fea56a",
   4745 => x"ffffff",
   4746 => x"ffffff",
   4747 => x"ffffff",
   4748 => x"ffffff",
   4749 => x"ffffff",
   4750 => x"ffffff",
   4751 => x"ffffff",
   4752 => x"ffffff",
   4753 => x"ffffff",
   4754 => x"ffffff",
   4755 => x"ffffff",
   4756 => x"ffffff",
   4757 => x"ffffff",
   4758 => x"ffffff",
   4759 => x"ffffff",
   4760 => x"ffffff",
   4761 => x"ffffff",
   4762 => x"ffffff",
   4763 => x"ffffff",
   4764 => x"ffffff",
   4765 => x"ffffff",
   4766 => x"ffffff",
   4767 => x"ffffff",
   4768 => x"ffffff",
   4769 => x"ffffff",
   4770 => x"ffffff",
   4771 => x"ffffff",
   4772 => x"ffffff",
   4773 => x"ffffff",
   4774 => x"ffffff",
   4775 => x"ffffff",
   4776 => x"ffffff",
   4777 => x"ffffff",
   4778 => x"ffffff",
   4779 => x"ffffff",
   4780 => x"ffffff",
   4781 => x"ffffff",
   4782 => x"ffffff",
   4783 => x"ffffff",
   4784 => x"ffffff",
   4785 => x"ffffff",
   4786 => x"ffffff",
   4787 => x"ffffff",
   4788 => x"ffffff",
   4789 => x"ffffff",
   4790 => x"ffffff",
   4791 => x"ffffff",
   4792 => x"ffffff",
   4793 => x"ffffff",
   4794 => x"ffffff",
   4795 => x"ffffff",
   4796 => x"ffffff",
   4797 => x"ffffff",
   4798 => x"ffffff",
   4799 => x"ffffff",
   4800 => x"ffffff",
   4801 => x"fff540",
   4802 => x"000abf",
   4803 => x"ffffff",
   4804 => x"ffffff",
   4805 => x"fff540",
   4806 => x"00057f",
   4807 => x"ffffff",
   4808 => x"ffffff",
   4809 => x"fffd70",
   4810 => x"c30c30",
   4811 => x"c30c30",
   4812 => x"c30c30",
   4813 => x"c30c30",
   4814 => x"c30c30",
   4815 => x"c30c30",
   4816 => x"c30c30",
   4817 => x"c30c30",
   4818 => x"c30c30",
   4819 => x"c30c30",
   4820 => x"c30c30",
   4821 => x"c30c30",
   4822 => x"c30c30",
   4823 => x"c30c30",
   4824 => x"c30c30",
   4825 => x"c30c30",
   4826 => x"c30c30",
   4827 => x"c30c30",
   4828 => x"c30c30",
   4829 => x"c30c30",
   4830 => x"c30c30",
   4831 => x"c2473c",
   4832 => x"f3cf3c",
   4833 => x"f3cf3c",
   4834 => x"f3cf3c",
   4835 => x"f3cf3c",
   4836 => x"f3cf2c",
   4837 => x"70c30c",
   4838 => x"30c30c",
   4839 => x"30c30c",
   4840 => x"30c30c",
   4841 => x"30c30c",
   4842 => x"30c30c",
   4843 => x"30c30c",
   4844 => x"30c30c",
   4845 => x"30c30c",
   4846 => x"30c30c",
   4847 => x"30c30c",
   4848 => x"30c30c",
   4849 => x"30c30c",
   4850 => x"30c30c",
   4851 => x"30c30c",
   4852 => x"30c30c",
   4853 => x"30c30c",
   4854 => x"30c30c",
   4855 => x"30c30c",
   4856 => x"30c30c",
   4857 => x"30c30c",
   4858 => x"30c31d",
   4859 => x"bbffff",
   4860 => x"ffffff",
   4861 => x"ffffff",
   4862 => x"a80000",
   4863 => x"00057f",
   4864 => x"ffffff",
   4865 => x"ffffff",
   4866 => x"fffa95",
   4867 => x"000015",
   4868 => x"ffffff",
   4869 => x"ffffff",
   4870 => x"ffffff",
   4871 => x"ffffff",
   4872 => x"ffffff",
   4873 => x"ffffff",
   4874 => x"ffffff",
   4875 => x"ffffff",
   4876 => x"ffffff",
   4877 => x"ffffff",
   4878 => x"ffffff",
   4879 => x"ffffff",
   4880 => x"ffffff",
   4881 => x"ffffff",
   4882 => x"ffffff",
   4883 => x"ffffff",
   4884 => x"ffffff",
   4885 => x"ffffff",
   4886 => x"ffffff",
   4887 => x"ffffff",
   4888 => x"ffffff",
   4889 => x"ffffff",
   4890 => x"ffffff",
   4891 => x"ffffff",
   4892 => x"ffffff",
   4893 => x"ffffff",
   4894 => x"ffffff",
   4895 => x"ffffff",
   4896 => x"ffffff",
   4897 => x"ffffff",
   4898 => x"ffffff",
   4899 => x"ffffff",
   4900 => x"ffffff",
   4901 => x"ffffff",
   4902 => x"ffffff",
   4903 => x"ffffff",
   4904 => x"a95abf",
   4905 => x"ffffff",
   4906 => x"ffffff",
   4907 => x"ffffff",
   4908 => x"ffffff",
   4909 => x"ffffff",
   4910 => x"ffffff",
   4911 => x"ffffff",
   4912 => x"ffffff",
   4913 => x"ffffff",
   4914 => x"ffffff",
   4915 => x"ffffff",
   4916 => x"ffffff",
   4917 => x"ffffff",
   4918 => x"ffffff",
   4919 => x"ffffff",
   4920 => x"ffffff",
   4921 => x"ffffff",
   4922 => x"ffffff",
   4923 => x"ffffff",
   4924 => x"ffffff",
   4925 => x"ffffff",
   4926 => x"ffffff",
   4927 => x"ffffff",
   4928 => x"ffffff",
   4929 => x"ffffff",
   4930 => x"ffffff",
   4931 => x"ffffff",
   4932 => x"ffffff",
   4933 => x"ffffff",
   4934 => x"ffffff",
   4935 => x"ffffff",
   4936 => x"ffffff",
   4937 => x"ffffff",
   4938 => x"ffffff",
   4939 => x"ffffff",
   4940 => x"ffffff",
   4941 => x"ffffff",
   4942 => x"ffffff",
   4943 => x"ffffff",
   4944 => x"ffffff",
   4945 => x"ffffff",
   4946 => x"ffffff",
   4947 => x"ffffff",
   4948 => x"ffffff",
   4949 => x"ffffff",
   4950 => x"ffffff",
   4951 => x"ffffff",
   4952 => x"ffffff",
   4953 => x"ffffff",
   4954 => x"ffffff",
   4955 => x"ffffff",
   4956 => x"ffffff",
   4957 => x"ffffff",
   4958 => x"ffffff",
   4959 => x"ffffff",
   4960 => x"ffffff",
   4961 => x"fff540",
   4962 => x"000abf",
   4963 => x"ffffff",
   4964 => x"ffffff",
   4965 => x"fffa80",
   4966 => x"00002a",
   4967 => x"ffffff",
   4968 => x"ffffff",
   4969 => x"eb5c30",
   4970 => x"c30c30",
   4971 => x"c30c30",
   4972 => x"c30c30",
   4973 => x"c30c30",
   4974 => x"c30c30",
   4975 => x"c30c30",
   4976 => x"c30c30",
   4977 => x"c30c30",
   4978 => x"c30c30",
   4979 => x"c30c30",
   4980 => x"c30c30",
   4981 => x"c30c30",
   4982 => x"c30c30",
   4983 => x"c30c30",
   4984 => x"c30c30",
   4985 => x"c30c30",
   4986 => x"c30c30",
   4987 => x"c30c30",
   4988 => x"c30c30",
   4989 => x"c30c30",
   4990 => x"c30c30",
   4991 => x"a2cf3c",
   4992 => x"f3cf3c",
   4993 => x"f3cf3c",
   4994 => x"f3cf3c",
   4995 => x"f3cf3c",
   4996 => x"f3cf3c",
   4997 => x"b1c30c",
   4998 => x"30c30c",
   4999 => x"30c30c",
   5000 => x"30c30c",
   5001 => x"30c30c",
   5002 => x"30c30c",
   5003 => x"30c30c",
   5004 => x"30c30c",
   5005 => x"30c30c",
   5006 => x"30c30c",
   5007 => x"30c30c",
   5008 => x"30c30c",
   5009 => x"30c30c",
   5010 => x"30c30c",
   5011 => x"30c30c",
   5012 => x"30c30c",
   5013 => x"30c30c",
   5014 => x"30c30c",
   5015 => x"30c30c",
   5016 => x"30c30c",
   5017 => x"30c30c",
   5018 => x"30c30c",
   5019 => x"31dfff",
   5020 => x"ffffff",
   5021 => x"ffffff",
   5022 => x"fea000",
   5023 => x"000015",
   5024 => x"56aaaa",
   5025 => x"aaaaaa",
   5026 => x"a95000",
   5027 => x"000015",
   5028 => x"ffffff",
   5029 => x"ffffff",
   5030 => x"ffffff",
   5031 => x"ffffff",
   5032 => x"ffffff",
   5033 => x"ffffff",
   5034 => x"ffffff",
   5035 => x"ffffff",
   5036 => x"ffffff",
   5037 => x"ffffff",
   5038 => x"ffffff",
   5039 => x"ffffff",
   5040 => x"ffffff",
   5041 => x"ffffff",
   5042 => x"ffffff",
   5043 => x"ffffff",
   5044 => x"ffffff",
   5045 => x"ffffff",
   5046 => x"ffffff",
   5047 => x"ffffff",
   5048 => x"ffffff",
   5049 => x"ffffff",
   5050 => x"ffffff",
   5051 => x"ffffff",
   5052 => x"ffffff",
   5053 => x"ffffff",
   5054 => x"ffffff",
   5055 => x"ffffff",
   5056 => x"ffffff",
   5057 => x"ffffff",
   5058 => x"ffffff",
   5059 => x"ffffff",
   5060 => x"ffffff",
   5061 => x"ffffff",
   5062 => x"ffffff",
   5063 => x"ffffea",
   5064 => x"56afff",
   5065 => x"ffffff",
   5066 => x"ffffff",
   5067 => x"ffffff",
   5068 => x"ffffff",
   5069 => x"ffffff",
   5070 => x"ffffff",
   5071 => x"ffffff",
   5072 => x"ffffff",
   5073 => x"ffffff",
   5074 => x"ffffff",
   5075 => x"ffffff",
   5076 => x"ffffff",
   5077 => x"ffffff",
   5078 => x"ffffff",
   5079 => x"ffffff",
   5080 => x"ffffff",
   5081 => x"ffffff",
   5082 => x"ffffff",
   5083 => x"ffffff",
   5084 => x"ffffff",
   5085 => x"ffffff",
   5086 => x"ffffff",
   5087 => x"ffffff",
   5088 => x"ffffff",
   5089 => x"ffffff",
   5090 => x"ffffff",
   5091 => x"ffffff",
   5092 => x"ffffff",
   5093 => x"ffffff",
   5094 => x"ffffff",
   5095 => x"ffffff",
   5096 => x"ffffff",
   5097 => x"ffffff",
   5098 => x"ffffff",
   5099 => x"ffffff",
   5100 => x"ffffff",
   5101 => x"ffffff",
   5102 => x"ffffff",
   5103 => x"ffffff",
   5104 => x"ffffff",
   5105 => x"ffffff",
   5106 => x"ffffff",
   5107 => x"ffffff",
   5108 => x"ffffff",
   5109 => x"ffffff",
   5110 => x"ffffff",
   5111 => x"ffffff",
   5112 => x"ffffff",
   5113 => x"ffffff",
   5114 => x"ffffff",
   5115 => x"ffffff",
   5116 => x"ffffff",
   5117 => x"ffffff",
   5118 => x"ffffff",
   5119 => x"ffffff",
   5120 => x"ffffff",
   5121 => x"fff540",
   5122 => x"000abf",
   5123 => x"ffffff",
   5124 => x"ffffff",
   5125 => x"ffffd5",
   5126 => x"000015",
   5127 => x"ffffff",
   5128 => x"fffffa",
   5129 => x"d70c30",
   5130 => x"c30c30",
   5131 => x"c30c30",
   5132 => x"c30c30",
   5133 => x"c30c30",
   5134 => x"c30c30",
   5135 => x"c30c30",
   5136 => x"c30c30",
   5137 => x"c30c30",
   5138 => x"c30c30",
   5139 => x"c30c30",
   5140 => x"c30c30",
   5141 => x"c30c30",
   5142 => x"c30c30",
   5143 => x"c30c30",
   5144 => x"c30c30",
   5145 => x"c30c30",
   5146 => x"c30c30",
   5147 => x"c30c30",
   5148 => x"c30c30",
   5149 => x"c30c30",
   5150 => x"c30918",
   5151 => x"b3cf3c",
   5152 => x"f3cf3c",
   5153 => x"f3cf3c",
   5154 => x"f3cf3c",
   5155 => x"f3cf3c",
   5156 => x"f3cf3c",
   5157 => x"f3cb0c",
   5158 => x"30c30c",
   5159 => x"30c30c",
   5160 => x"30c30c",
   5161 => x"30c30c",
   5162 => x"30c30c",
   5163 => x"30c30c",
   5164 => x"30c30c",
   5165 => x"30c30c",
   5166 => x"30c30c",
   5167 => x"30c30c",
   5168 => x"30c30c",
   5169 => x"30c30c",
   5170 => x"30c30c",
   5171 => x"30c30c",
   5172 => x"30c30c",
   5173 => x"30c30c",
   5174 => x"30c30c",
   5175 => x"30c30c",
   5176 => x"30c30c",
   5177 => x"30c30c",
   5178 => x"30c30c",
   5179 => x"30c77f",
   5180 => x"ffffff",
   5181 => x"ffffff",
   5182 => x"fffa95",
   5183 => x"000000",
   5184 => x"000000",
   5185 => x"555000",
   5186 => x"000000",
   5187 => x"00056a",
   5188 => x"ffffff",
   5189 => x"ffffff",
   5190 => x"ffffff",
   5191 => x"ffffff",
   5192 => x"ffffff",
   5193 => x"ffffff",
   5194 => x"ffffff",
   5195 => x"ffffff",
   5196 => x"ffffff",
   5197 => x"ffffff",
   5198 => x"ffffff",
   5199 => x"ffffff",
   5200 => x"ffffff",
   5201 => x"ffffff",
   5202 => x"ffffff",
   5203 => x"ffffff",
   5204 => x"ffffff",
   5205 => x"ffffff",
   5206 => x"ffffff",
   5207 => x"ffffff",
   5208 => x"ffffff",
   5209 => x"ffffff",
   5210 => x"ffffff",
   5211 => x"ffffff",
   5212 => x"ffffff",
   5213 => x"ffffff",
   5214 => x"ffffff",
   5215 => x"ffffff",
   5216 => x"ffffff",
   5217 => x"ffffff",
   5218 => x"ffffff",
   5219 => x"ffffff",
   5220 => x"ffffff",
   5221 => x"ffffff",
   5222 => x"ffffff",
   5223 => x"fffa95",
   5224 => x"abffff",
   5225 => x"ffffff",
   5226 => x"ffffff",
   5227 => x"ffffff",
   5228 => x"ffffff",
   5229 => x"ffffff",
   5230 => x"ffffff",
   5231 => x"ffffff",
   5232 => x"ffffff",
   5233 => x"ffffff",
   5234 => x"ffffff",
   5235 => x"ffffff",
   5236 => x"ffffff",
   5237 => x"ffffff",
   5238 => x"ffffff",
   5239 => x"ffffff",
   5240 => x"ffffff",
   5241 => x"ffffff",
   5242 => x"ffffff",
   5243 => x"ffffff",
   5244 => x"ffffff",
   5245 => x"ffffff",
   5246 => x"ffffff",
   5247 => x"ffffff",
   5248 => x"ffffff",
   5249 => x"ffffff",
   5250 => x"ffffff",
   5251 => x"ffffff",
   5252 => x"ffffff",
   5253 => x"ffffff",
   5254 => x"ffffff",
   5255 => x"ffffff",
   5256 => x"ffffff",
   5257 => x"ffffff",
   5258 => x"ffffff",
   5259 => x"ffffff",
   5260 => x"ffffff",
   5261 => x"ffffff",
   5262 => x"ffffff",
   5263 => x"ffffff",
   5264 => x"ffffff",
   5265 => x"ffffff",
   5266 => x"ffffff",
   5267 => x"ffffff",
   5268 => x"ffffff",
   5269 => x"ffffff",
   5270 => x"ffffff",
   5271 => x"ffffff",
   5272 => x"ffffff",
   5273 => x"ffffff",
   5274 => x"ffffff",
   5275 => x"ffffff",
   5276 => x"ffffff",
   5277 => x"ffffff",
   5278 => x"ffffff",
   5279 => x"ffffff",
   5280 => x"ffffff",
   5281 => x"fff540",
   5282 => x"000abf",
   5283 => x"ffffff",
   5284 => x"ffffff",
   5285 => x"ffffea",
   5286 => x"000000",
   5287 => x"abffff",
   5288 => x"fffeb0",
   5289 => x"c30c30",
   5290 => x"c30c30",
   5291 => x"c30c30",
   5292 => x"c30c30",
   5293 => x"c30c30",
   5294 => x"c30c30",
   5295 => x"c30c30",
   5296 => x"c30c30",
   5297 => x"c30c30",
   5298 => x"c30c30",
   5299 => x"c30c30",
   5300 => x"c30c30",
   5301 => x"c30c30",
   5302 => x"c30c30",
   5303 => x"c30c30",
   5304 => x"c30c30",
   5305 => x"c30c30",
   5306 => x"c30c30",
   5307 => x"c30c30",
   5308 => x"c30c30",
   5309 => x"c30c30",
   5310 => x"c24a2c",
   5311 => x"f3cf3c",
   5312 => x"f3cf3c",
   5313 => x"f3cf3c",
   5314 => x"f3cf3c",
   5315 => x"f3cf3c",
   5316 => x"f3cf3c",
   5317 => x"f3cf2c",
   5318 => x"70c30c",
   5319 => x"30c30c",
   5320 => x"30c30c",
   5321 => x"30c30c",
   5322 => x"30c30c",
   5323 => x"30c30c",
   5324 => x"30c30c",
   5325 => x"30c30c",
   5326 => x"30c30c",
   5327 => x"30c30c",
   5328 => x"30c30c",
   5329 => x"30c30c",
   5330 => x"30c30c",
   5331 => x"30c30c",
   5332 => x"30c30c",
   5333 => x"30c30c",
   5334 => x"30c30c",
   5335 => x"30c30c",
   5336 => x"30c30c",
   5337 => x"30c30c",
   5338 => x"30c30c",
   5339 => x"30c31d",
   5340 => x"bbffff",
   5341 => x"ffffff",
   5342 => x"ffffea",
   5343 => x"a95000",
   5344 => x"000000",
   5345 => x"000000",
   5346 => x"000000",
   5347 => x"56afff",
   5348 => x"ffffff",
   5349 => x"ffffff",
   5350 => x"ffffff",
   5351 => x"ffffff",
   5352 => x"ffffff",
   5353 => x"ffffff",
   5354 => x"ffffff",
   5355 => x"ffffff",
   5356 => x"ffffff",
   5357 => x"ffffff",
   5358 => x"ffffff",
   5359 => x"ffffff",
   5360 => x"ffffff",
   5361 => x"ffffff",
   5362 => x"ffffff",
   5363 => x"ffffff",
   5364 => x"ffffff",
   5365 => x"ffffff",
   5366 => x"ffffff",
   5367 => x"ffffff",
   5368 => x"ffffff",
   5369 => x"ffffff",
   5370 => x"ffffff",
   5371 => x"ffffff",
   5372 => x"ffffff",
   5373 => x"ffffff",
   5374 => x"ffffff",
   5375 => x"ffffff",
   5376 => x"ffffff",
   5377 => x"ffffff",
   5378 => x"ffffff",
   5379 => x"ffffff",
   5380 => x"ffffff",
   5381 => x"ffffff",
   5382 => x"ffffff",
   5383 => x"fea56a",
   5384 => x"ffffff",
   5385 => x"ffffff",
   5386 => x"ffffff",
   5387 => x"ffffff",
   5388 => x"ffffff",
   5389 => x"ffffff",
   5390 => x"ffffff",
   5391 => x"ffffff",
   5392 => x"ffffff",
   5393 => x"ffffff",
   5394 => x"ffffff",
   5395 => x"ffffff",
   5396 => x"ffffff",
   5397 => x"ffffff",
   5398 => x"ffffff",
   5399 => x"ffffff",
   5400 => x"ffffff",
   5401 => x"ffffff",
   5402 => x"ffffff",
   5403 => x"ffffff",
   5404 => x"ffffff",
   5405 => x"ffffff",
   5406 => x"ffffff",
   5407 => x"ffffff",
   5408 => x"ffffff",
   5409 => x"ffffff",
   5410 => x"ffffff",
   5411 => x"ffffff",
   5412 => x"ffffff",
   5413 => x"ffffff",
   5414 => x"ffffff",
   5415 => x"ffffff",
   5416 => x"ffffff",
   5417 => x"ffffff",
   5418 => x"ffffff",
   5419 => x"ffffff",
   5420 => x"ffffff",
   5421 => x"ffffff",
   5422 => x"ffffff",
   5423 => x"ffffff",
   5424 => x"ffffff",
   5425 => x"ffffff",
   5426 => x"ffffff",
   5427 => x"ffffff",
   5428 => x"ffffff",
   5429 => x"ffffff",
   5430 => x"ffffff",
   5431 => x"ffffff",
   5432 => x"ffffff",
   5433 => x"ffffff",
   5434 => x"ffffff",
   5435 => x"ffffff",
   5436 => x"ffffff",
   5437 => x"ffffff",
   5438 => x"ffffff",
   5439 => x"ffffff",
   5440 => x"ffffff",
   5441 => x"fff540",
   5442 => x"000abf",
   5443 => x"ffffff",
   5444 => x"ffffff",
   5445 => x"ffffff",
   5446 => x"540000",
   5447 => x"57ffff",
   5448 => x"ff5c30",
   5449 => x"c30c30",
   5450 => x"c30c30",
   5451 => x"c30c30",
   5452 => x"c30c30",
   5453 => x"c30c30",
   5454 => x"c30c30",
   5455 => x"c30c30",
   5456 => x"c30c30",
   5457 => x"c30c30",
   5458 => x"c30c30",
   5459 => x"c30c30",
   5460 => x"c30c30",
   5461 => x"c30c30",
   5462 => x"c30c30",
   5463 => x"c30c30",
   5464 => x"c30c30",
   5465 => x"c30c30",
   5466 => x"c30c30",
   5467 => x"c30c30",
   5468 => x"c30c30",
   5469 => x"c30c30",
   5470 => x"92cf3c",
   5471 => x"f3cf3c",
   5472 => x"f3cf3c",
   5473 => x"f3cf3c",
   5474 => x"f3cf3c",
   5475 => x"f3cf3c",
   5476 => x"f3cf3c",
   5477 => x"f3cf3c",
   5478 => x"b1c30c",
   5479 => x"30c30c",
   5480 => x"30c30c",
   5481 => x"30c30c",
   5482 => x"30c30c",
   5483 => x"30c30c",
   5484 => x"30c30c",
   5485 => x"30c30c",
   5486 => x"30c30c",
   5487 => x"30c30c",
   5488 => x"30c30c",
   5489 => x"30c30c",
   5490 => x"30c30c",
   5491 => x"30c30c",
   5492 => x"30c30c",
   5493 => x"30c30c",
   5494 => x"30c30c",
   5495 => x"30c30c",
   5496 => x"30c30c",
   5497 => x"30c30c",
   5498 => x"30c30c",
   5499 => x"30c30c",
   5500 => x"76efff",
   5501 => x"ffffff",
   5502 => x"ffffff",
   5503 => x"feaa95",
   5504 => x"540000",
   5505 => x"000000",
   5506 => x"555aaa",
   5507 => x"ffffff",
   5508 => x"ffffff",
   5509 => x"ffffff",
   5510 => x"ffffff",
   5511 => x"ffffff",
   5512 => x"ffffff",
   5513 => x"ffffff",
   5514 => x"ffffff",
   5515 => x"ffffff",
   5516 => x"ffffff",
   5517 => x"ffffff",
   5518 => x"ffffff",
   5519 => x"ffffff",
   5520 => x"ffffff",
   5521 => x"ffffff",
   5522 => x"ffffff",
   5523 => x"ffffff",
   5524 => x"ffffff",
   5525 => x"ffffff",
   5526 => x"ffffff",
   5527 => x"ffffff",
   5528 => x"ffffff",
   5529 => x"ffffff",
   5530 => x"ffffff",
   5531 => x"ffffff",
   5532 => x"ffffff",
   5533 => x"ffffff",
   5534 => x"ffffff",
   5535 => x"ffffff",
   5536 => x"ffffff",
   5537 => x"ffffff",
   5538 => x"ffffff",
   5539 => x"ffffff",
   5540 => x"ffffff",
   5541 => x"ffffff",
   5542 => x"ffffff",
   5543 => x"a95abf",
   5544 => x"ffffff",
   5545 => x"ffffff",
   5546 => x"ffffff",
   5547 => x"ffffff",
   5548 => x"ffffff",
   5549 => x"ffffff",
   5550 => x"ffffff",
   5551 => x"ffffff",
   5552 => x"ffffff",
   5553 => x"ffffff",
   5554 => x"ffffff",
   5555 => x"ffffff",
   5556 => x"ffffff",
   5557 => x"ffffff",
   5558 => x"ffffff",
   5559 => x"ffffff",
   5560 => x"ffffff",
   5561 => x"ffffff",
   5562 => x"ffffff",
   5563 => x"ffffff",
   5564 => x"ffffff",
   5565 => x"ffffff",
   5566 => x"ffffff",
   5567 => x"ffffff",
   5568 => x"ffffff",
   5569 => x"ffffff",
   5570 => x"ffffff",
   5571 => x"ffffff",
   5572 => x"ffffff",
   5573 => x"ffffff",
   5574 => x"ffffff",
   5575 => x"ffffff",
   5576 => x"ffffff",
   5577 => x"ffffff",
   5578 => x"ffffff",
   5579 => x"ffffff",
   5580 => x"ffffff",
   5581 => x"ffffff",
   5582 => x"ffffff",
   5583 => x"ffffff",
   5584 => x"ffffff",
   5585 => x"ffffff",
   5586 => x"ffffff",
   5587 => x"ffffff",
   5588 => x"ffffff",
   5589 => x"ffffff",
   5590 => x"ffffff",
   5591 => x"ffffff",
   5592 => x"ffffff",
   5593 => x"ffffff",
   5594 => x"ffffff",
   5595 => x"ffffff",
   5596 => x"ffffff",
   5597 => x"ffffff",
   5598 => x"ffffff",
   5599 => x"ffffff",
   5600 => x"ffffff",
   5601 => x"fff540",
   5602 => x"000abf",
   5603 => x"ffffff",
   5604 => x"ffffff",
   5605 => x"ffffff",
   5606 => x"a80000",
   5607 => x"02afff",
   5608 => x"d70c30",
   5609 => x"c30c30",
   5610 => x"c30c30",
   5611 => x"c30c30",
   5612 => x"c30c30",
   5613 => x"c30c30",
   5614 => x"c30c30",
   5615 => x"c30c30",
   5616 => x"c30c30",
   5617 => x"c30c30",
   5618 => x"c30c30",
   5619 => x"c30c30",
   5620 => x"c30c30",
   5621 => x"c30c30",
   5622 => x"c30c30",
   5623 => x"c30c30",
   5624 => x"c30c30",
   5625 => x"c30c30",
   5626 => x"c30c30",
   5627 => x"c30c30",
   5628 => x"c30c30",
   5629 => x"c30c24",
   5630 => x"b3cf3c",
   5631 => x"f3cf3c",
   5632 => x"f3cf3c",
   5633 => x"f3cf3c",
   5634 => x"f3cf3c",
   5635 => x"f3cf3c",
   5636 => x"f3cf3c",
   5637 => x"f3cf3c",
   5638 => x"f2c70c",
   5639 => x"30c30c",
   5640 => x"30c30c",
   5641 => x"30c30c",
   5642 => x"30c30c",
   5643 => x"30c30c",
   5644 => x"30c30c",
   5645 => x"30c30c",
   5646 => x"30c30c",
   5647 => x"30c30c",
   5648 => x"30c30c",
   5649 => x"30c30c",
   5650 => x"30c30c",
   5651 => x"30c30c",
   5652 => x"30c30c",
   5653 => x"30c30c",
   5654 => x"30c30c",
   5655 => x"30c30c",
   5656 => x"30c30c",
   5657 => x"30c30c",
   5658 => x"30c30c",
   5659 => x"30c30c",
   5660 => x"31dbbf",
   5661 => x"ffffff",
   5662 => x"ffffff",
   5663 => x"ffffff",
   5664 => x"aaaaaa",
   5665 => x"aaaaaa",
   5666 => x"abffff",
   5667 => x"ffffff",
   5668 => x"ffffff",
   5669 => x"ffffff",
   5670 => x"ffffff",
   5671 => x"ffffff",
   5672 => x"ffffff",
   5673 => x"ffffff",
   5674 => x"ffffff",
   5675 => x"ffffff",
   5676 => x"ffffff",
   5677 => x"ffffff",
   5678 => x"ffffff",
   5679 => x"ffffff",
   5680 => x"ffffff",
   5681 => x"ffffff",
   5682 => x"ffffff",
   5683 => x"ffffff",
   5684 => x"ffffff",
   5685 => x"ffffff",
   5686 => x"ffffff",
   5687 => x"ffffff",
   5688 => x"ffffff",
   5689 => x"ffffff",
   5690 => x"ffffff",
   5691 => x"ffffff",
   5692 => x"ffffff",
   5693 => x"ffffff",
   5694 => x"ffffff",
   5695 => x"ffffff",
   5696 => x"ffffff",
   5697 => x"ffffff",
   5698 => x"ffffff",
   5699 => x"ffffff",
   5700 => x"ffffff",
   5701 => x"ffffff",
   5702 => x"ffffea",
   5703 => x"56afff",
   5704 => x"ffffff",
   5705 => x"ffffff",
   5706 => x"ffffff",
   5707 => x"ffffff",
   5708 => x"ffffff",
   5709 => x"ffffff",
   5710 => x"ffffff",
   5711 => x"ffffff",
   5712 => x"ffffff",
   5713 => x"ffffff",
   5714 => x"ffffff",
   5715 => x"ffffff",
   5716 => x"ffffff",
   5717 => x"ffffff",
   5718 => x"ffffff",
   5719 => x"ffffff",
   5720 => x"ffffff",
   5721 => x"ffffff",
   5722 => x"ffffff",
   5723 => x"ffffff",
   5724 => x"ffffff",
   5725 => x"ffffff",
   5726 => x"ffffff",
   5727 => x"ffffff",
   5728 => x"ffffff",
   5729 => x"ffffff",
   5730 => x"ffffff",
   5731 => x"ffffff",
   5732 => x"ffffff",
   5733 => x"ffffff",
   5734 => x"ffffff",
   5735 => x"ffffff",
   5736 => x"ffffff",
   5737 => x"ffffff",
   5738 => x"ffffff",
   5739 => x"ffffff",
   5740 => x"ffffff",
   5741 => x"ffffff",
   5742 => x"ffffff",
   5743 => x"ffffff",
   5744 => x"ffffff",
   5745 => x"ffffff",
   5746 => x"ffffff",
   5747 => x"ffffff",
   5748 => x"ffffff",
   5749 => x"ffffff",
   5750 => x"ffffff",
   5751 => x"ffffff",
   5752 => x"ffffff",
   5753 => x"ffffff",
   5754 => x"ffffff",
   5755 => x"ffffff",
   5756 => x"ffffff",
   5757 => x"ffffff",
   5758 => x"ffffff",
   5759 => x"ffffff",
   5760 => x"ffffff",
   5761 => x"fffa95",
   5762 => x"56afff",
   5763 => x"ffffff",
   5764 => x"ffffff",
   5765 => x"ffffff",
   5766 => x"fea555",
   5767 => x"56aff5",
   5768 => x"c30c30",
   5769 => x"c30c30",
   5770 => x"c30c30",
   5771 => x"c30c30",
   5772 => x"c30c30",
   5773 => x"c30c30",
   5774 => x"c30c30",
   5775 => x"c30c30",
   5776 => x"c30c30",
   5777 => x"c30c30",
   5778 => x"c30c30",
   5779 => x"c30c30",
   5780 => x"c30c30",
   5781 => x"c30c30",
   5782 => x"c30c30",
   5783 => x"c30c30",
   5784 => x"c30c30",
   5785 => x"c30c30",
   5786 => x"c30c30",
   5787 => x"c30c30",
   5788 => x"c30c30",
   5789 => x"c30a2c",
   5790 => x"f3cf3c",
   5791 => x"f3cf3c",
   5792 => x"f3cf3c",
   5793 => x"f3cf3c",
   5794 => x"f3cf3c",
   5795 => x"f3cf3c",
   5796 => x"f3cf3c",
   5797 => x"f3cf3c",
   5798 => x"f3cb1c",
   5799 => x"30c30c",
   5800 => x"30c30c",
   5801 => x"30c30c",
   5802 => x"30c30c",
   5803 => x"30c30c",
   5804 => x"30c30c",
   5805 => x"30c30c",
   5806 => x"30c30c",
   5807 => x"30c30c",
   5808 => x"30c30c",
   5809 => x"30c30c",
   5810 => x"30c30c",
   5811 => x"30c30c",
   5812 => x"30c30c",
   5813 => x"30c30c",
   5814 => x"30c30c",
   5815 => x"30c30c",
   5816 => x"30c30c",
   5817 => x"30c30c",
   5818 => x"30c30c",
   5819 => x"30c30c",
   5820 => x"30c32e",
   5821 => x"ffffff",
   5822 => x"ffffff",
   5823 => x"ffffff",
   5824 => x"ffffff",
   5825 => x"ffffff",
   5826 => x"ffffff",
   5827 => x"ffffff",
   5828 => x"ffffff",
   5829 => x"ffffff",
   5830 => x"ffffff",
   5831 => x"ffffff",
   5832 => x"ffffff",
   5833 => x"ffffff",
   5834 => x"ffffff",
   5835 => x"ffffff",
   5836 => x"ffffff",
   5837 => x"ffffff",
   5838 => x"ffffff",
   5839 => x"ffffff",
   5840 => x"ffffff",
   5841 => x"ffffff",
   5842 => x"ffffff",
   5843 => x"ffffff",
   5844 => x"ffffff",
   5845 => x"ffffff",
   5846 => x"ffffff",
   5847 => x"ffffff",
   5848 => x"ffffff",
   5849 => x"ffffff",
   5850 => x"ffffff",
   5851 => x"ffffff",
   5852 => x"ffffff",
   5853 => x"ffffff",
   5854 => x"ffffff",
   5855 => x"ffffff",
   5856 => x"ffffff",
   5857 => x"ffffff",
   5858 => x"ffffff",
   5859 => x"ffffff",
   5860 => x"ffffff",
   5861 => x"ffffff",
   5862 => x"fffa95",
   5863 => x"abffff",
   5864 => x"ffffff",
   5865 => x"ffffff",
   5866 => x"ffffff",
   5867 => x"ffffff",
   5868 => x"ffffff",
   5869 => x"ffffff",
   5870 => x"ffffff",
   5871 => x"ffffff",
   5872 => x"ffffff",
   5873 => x"ffffff",
   5874 => x"ffffff",
   5875 => x"ffffff",
   5876 => x"ffffff",
   5877 => x"ffffff",
   5878 => x"ffffff",
   5879 => x"ffffff",
   5880 => x"ffffff",
   5881 => x"ffffff",
   5882 => x"ffffff",
   5883 => x"ffffff",
   5884 => x"ffffff",
   5885 => x"ffffff",
   5886 => x"ffffff",
   5887 => x"ffffff",
   5888 => x"ffffff",
   5889 => x"ffffff",
   5890 => x"ffffff",
   5891 => x"ffffff",
   5892 => x"ffffff",
   5893 => x"ffffff",
   5894 => x"ffffff",
   5895 => x"ffffff",
   5896 => x"ffffff",
   5897 => x"ffffff",
   5898 => x"ffffff",
   5899 => x"ffffff",
   5900 => x"ffffff",
   5901 => x"ffffff",
   5902 => x"ffffff",
   5903 => x"ffffff",
   5904 => x"ffffff",
   5905 => x"ffffff",
   5906 => x"ffffff",
   5907 => x"ffffff",
   5908 => x"ffffff",
   5909 => x"ffffff",
   5910 => x"ffffff",
   5911 => x"ffffff",
   5912 => x"ffffff",
   5913 => x"ffffff",
   5914 => x"ffffff",
   5915 => x"ffffff",
   5916 => x"ffffff",
   5917 => x"ffffff",
   5918 => x"ffffff",
   5919 => x"ffffff",
   5920 => x"ffffff",
   5921 => x"ffffff",
   5922 => x"ffffff",
   5923 => x"ffffff",
   5924 => x"ffffff",
   5925 => x"ffffff",
   5926 => x"ffffff",
   5927 => x"ffad70",
   5928 => x"c30c30",
   5929 => x"c30c30",
   5930 => x"c30c30",
   5931 => x"c30c30",
   5932 => x"c30c30",
   5933 => x"c30c30",
   5934 => x"c30c30",
   5935 => x"c30c30",
   5936 => x"c30c30",
   5937 => x"c30c30",
   5938 => x"c30c30",
   5939 => x"c30c30",
   5940 => x"c30c30",
   5941 => x"c30c30",
   5942 => x"c30c30",
   5943 => x"c30c30",
   5944 => x"c30c30",
   5945 => x"c30c30",
   5946 => x"c30c30",
   5947 => x"c30c30",
   5948 => x"c30c30",
   5949 => x"c28b3c",
   5950 => x"f3cf3c",
   5951 => x"f3cf3c",
   5952 => x"f3cf3c",
   5953 => x"f3cf3c",
   5954 => x"f3cf3c",
   5955 => x"f3cf3c",
   5956 => x"f3cf3c",
   5957 => x"f3cf3c",
   5958 => x"f3cf3c",
   5959 => x"70c30c",
   5960 => x"30c30c",
   5961 => x"30c30c",
   5962 => x"30c30c",
   5963 => x"30c30c",
   5964 => x"30c30c",
   5965 => x"30c30c",
   5966 => x"30c30c",
   5967 => x"30c30c",
   5968 => x"30c30c",
   5969 => x"30c30c",
   5970 => x"30c30c",
   5971 => x"30c30c",
   5972 => x"30c30c",
   5973 => x"30c30c",
   5974 => x"30c30c",
   5975 => x"30c30c",
   5976 => x"30c30c",
   5977 => x"30c30c",
   5978 => x"30c30c",
   5979 => x"30c30c",
   5980 => x"30c30c",
   5981 => x"bbffff",
   5982 => x"ffffff",
   5983 => x"ffffff",
   5984 => x"ffffff",
   5985 => x"ffffff",
   5986 => x"ffffff",
   5987 => x"ffffff",
   5988 => x"ffffff",
   5989 => x"ffffff",
   5990 => x"ffffff",
   5991 => x"ffffff",
   5992 => x"ffffff",
   5993 => x"ffffff",
   5994 => x"ffffff",
   5995 => x"ffffff",
   5996 => x"ffffff",
   5997 => x"ffffff",
   5998 => x"ffffff",
   5999 => x"ffffff",
   6000 => x"ffffff",
   6001 => x"ffffff",
   6002 => x"ffffff",
   6003 => x"ffffff",
   6004 => x"ffffff",
   6005 => x"ffffff",
   6006 => x"ffffff",
   6007 => x"ffffff",
   6008 => x"ffffff",
   6009 => x"ffffff",
   6010 => x"ffffff",
   6011 => x"ffffff",
   6012 => x"ffffff",
   6013 => x"ffffff",
   6014 => x"ffffff",
   6015 => x"ffffff",
   6016 => x"ffffff",
   6017 => x"ffffff",
   6018 => x"ffffff",
   6019 => x"ffffff",
   6020 => x"ffffff",
   6021 => x"ffffff",
   6022 => x"fea56a",
   6023 => x"ffffff",
   6024 => x"ffffff",
   6025 => x"ffffff",
   6026 => x"ffffff",
   6027 => x"ffffff",
   6028 => x"ffffff",
   6029 => x"ffffff",
   6030 => x"ffffff",
   6031 => x"ffffff",
   6032 => x"ffffff",
   6033 => x"ffffff",
   6034 => x"ffffff",
   6035 => x"ffffff",
   6036 => x"ffffff",
   6037 => x"ffffff",
   6038 => x"ffffff",
   6039 => x"ffffff",
   6040 => x"ffffff",
   6041 => x"ffffff",
   6042 => x"ffffff",
   6043 => x"ffffff",
   6044 => x"ffffff",
   6045 => x"ffffff",
   6046 => x"ffffff",
   6047 => x"ffffff",
   6048 => x"ffffff",
   6049 => x"ffffff",
   6050 => x"ffffff",
   6051 => x"ffffff",
   6052 => x"ffffff",
   6053 => x"ffffff",
   6054 => x"ffffff",
   6055 => x"ffffff",
   6056 => x"ffffff",
   6057 => x"ffffff",
   6058 => x"ffffff",
   6059 => x"ffffff",
   6060 => x"ffffff",
   6061 => x"ffffff",
   6062 => x"ffffff",
   6063 => x"ffffff",
   6064 => x"ffffff",
   6065 => x"ffffff",
   6066 => x"ffffff",
   6067 => x"ffffff",
   6068 => x"ffffff",
   6069 => x"ffffff",
   6070 => x"ffffff",
   6071 => x"ffffff",
   6072 => x"ffffff",
   6073 => x"ffffff",
   6074 => x"ffffff",
   6075 => x"ffffff",
   6076 => x"ffffff",
   6077 => x"ffffff",
   6078 => x"ffffff",
   6079 => x"ffffff",
   6080 => x"ffffff",
   6081 => x"ffffff",
   6082 => x"ffffff",
   6083 => x"ffffff",
   6084 => x"ffffff",
   6085 => x"ffffff",
   6086 => x"ffffff",
   6087 => x"eb5c30",
   6088 => x"c30c30",
   6089 => x"c30c30",
   6090 => x"c30c30",
   6091 => x"c30c30",
   6092 => x"c30c30",
   6093 => x"c30c30",
   6094 => x"c30c30",
   6095 => x"c30c30",
   6096 => x"c30c30",
   6097 => x"c30c30",
   6098 => x"c30c30",
   6099 => x"c30c30",
   6100 => x"c30c30",
   6101 => x"c30c30",
   6102 => x"c30c30",
   6103 => x"c30c30",
   6104 => x"c30c30",
   6105 => x"c30c30",
   6106 => x"c30c30",
   6107 => x"c30c30",
   6108 => x"c30c24",
   6109 => x"a2cf3c",
   6110 => x"f3cf3c",
   6111 => x"f3cf3c",
   6112 => x"f3cf3c",
   6113 => x"f3cf3c",
   6114 => x"f3cf3c",
   6115 => x"f3cf3c",
   6116 => x"f3cf3c",
   6117 => x"f3cf3c",
   6118 => x"f3cf3c",
   6119 => x"f1c30c",
   6120 => x"30c30c",
   6121 => x"30c30c",
   6122 => x"30c30c",
   6123 => x"30c30c",
   6124 => x"30c30c",
   6125 => x"30c30c",
   6126 => x"30c30c",
   6127 => x"30c30c",
   6128 => x"30c30c",
   6129 => x"30c30c",
   6130 => x"30c30c",
   6131 => x"30c30c",
   6132 => x"30c30c",
   6133 => x"30c30c",
   6134 => x"30c30c",
   6135 => x"30c30c",
   6136 => x"30c30c",
   6137 => x"30c30c",
   6138 => x"30c30c",
   6139 => x"30c30c",
   6140 => x"30c30c",
   6141 => x"32efff",
   6142 => x"ffffff",
   6143 => x"ffffff",
   6144 => x"ffffff",
   6145 => x"ffffff",
   6146 => x"ffffff",
   6147 => x"ffffff",
   6148 => x"ffffff",
   6149 => x"ffffff",
   6150 => x"ffffff",
   6151 => x"ffffff",
   6152 => x"ffffff",
   6153 => x"ffffff",
   6154 => x"ffffff",
   6155 => x"ffffff",
   6156 => x"ffffff",
   6157 => x"ffffff",
   6158 => x"ffffff",
   6159 => x"ffffff",
   6160 => x"ffffff",
   6161 => x"ffffff",
   6162 => x"ffffff",
   6163 => x"ffffff",
   6164 => x"ffffff",
   6165 => x"ffffff",
   6166 => x"ffffff",
   6167 => x"ffffff",
   6168 => x"ffffff",
   6169 => x"ffffff",
   6170 => x"ffffff",
   6171 => x"ffffff",
   6172 => x"ffffff",
   6173 => x"ffffff",
   6174 => x"ffffff",
   6175 => x"ffffff",
   6176 => x"ffffff",
   6177 => x"ffffff",
   6178 => x"ffffff",
   6179 => x"ffffff",
   6180 => x"ffffff",
   6181 => x"ffffff",
   6182 => x"a95abf",
   6183 => x"ffffff",
   6184 => x"ffffff",
   6185 => x"ffffff",
   6186 => x"ffffff",
   6187 => x"ffffff",
   6188 => x"ffffff",
   6189 => x"ffffff",
   6190 => x"ffffff",
   6191 => x"ffffff",
   6192 => x"ffffff",
   6193 => x"ffffff",
   6194 => x"ffffff",
   6195 => x"ffffff",
   6196 => x"ffffff",
   6197 => x"ffffff",
   6198 => x"ffffff",
   6199 => x"ffffff",
   6200 => x"ffffff",
   6201 => x"ffffff",
   6202 => x"ffffff",
   6203 => x"ffffff",
   6204 => x"ffffff",
   6205 => x"ffffff",
   6206 => x"ffffff",
   6207 => x"ffffff",
   6208 => x"ffffff",
   6209 => x"ffffff",
   6210 => x"ffffff",
   6211 => x"ffffff",
   6212 => x"ffffff",
   6213 => x"ffffff",
   6214 => x"ffffff",
   6215 => x"ffffff",
   6216 => x"ffffff",
   6217 => x"ffffff",
   6218 => x"ffffff",
   6219 => x"ffffff",
   6220 => x"ffffff",
   6221 => x"ffffff",
   6222 => x"ffffff",
   6223 => x"ffffff",
   6224 => x"ffffff",
   6225 => x"ffffff",
   6226 => x"ffffff",
   6227 => x"ffffff",
   6228 => x"ffffff",
   6229 => x"ffffff",
   6230 => x"ffffff",
   6231 => x"ffffff",
   6232 => x"ffffff",
   6233 => x"ffffff",
   6234 => x"ffffff",
   6235 => x"ffffff",
   6236 => x"ffffff",
   6237 => x"ffffff",
   6238 => x"ffffff",
   6239 => x"ffffff",
   6240 => x"ffffff",
   6241 => x"ffffff",
   6242 => x"ffffff",
   6243 => x"ffffff",
   6244 => x"ffffff",
   6245 => x"ffffff",
   6246 => x"fffffa",
   6247 => x"d70c30",
   6248 => x"c30c30",
   6249 => x"c30c30",
   6250 => x"c30c30",
   6251 => x"c30c30",
   6252 => x"c30c30",
   6253 => x"c30c30",
   6254 => x"c30c30",
   6255 => x"c30c30",
   6256 => x"c30c30",
   6257 => x"c30c30",
   6258 => x"c30c30",
   6259 => x"c30c30",
   6260 => x"c30c30",
   6261 => x"c30c30",
   6262 => x"c30c30",
   6263 => x"c30c30",
   6264 => x"c30c30",
   6265 => x"c30c30",
   6266 => x"c30c30",
   6267 => x"c30c30",
   6268 => x"c30828",
   6269 => x"b3cf3c",
   6270 => x"f3cf3c",
   6271 => x"f3cf3c",
   6272 => x"f3cf3c",
   6273 => x"f3cf3c",
   6274 => x"f3cf3c",
   6275 => x"f3cf3c",
   6276 => x"f3cf3c",
   6277 => x"f3cf3c",
   6278 => x"f3cf3c",
   6279 => x"f3cb0c",
   6280 => x"30c30c",
   6281 => x"30c30c",
   6282 => x"30c30c",
   6283 => x"30c30c",
   6284 => x"30c30c",
   6285 => x"30c30c",
   6286 => x"30c30c",
   6287 => x"30c30c",
   6288 => x"30c30c",
   6289 => x"30c30c",
   6290 => x"30c30c",
   6291 => x"30c30c",
   6292 => x"30c30c",
   6293 => x"30c30c",
   6294 => x"30c30c",
   6295 => x"30c30c",
   6296 => x"30c30c",
   6297 => x"30c30c",
   6298 => x"30c30c",
   6299 => x"30c30c",
   6300 => x"30c30c",
   6301 => x"30c77f",
   6302 => x"ffffff",
   6303 => x"ffffff",
   6304 => x"ffffff",
   6305 => x"ffffff",
   6306 => x"ffffff",
   6307 => x"ffffff",
   6308 => x"ffffff",
   6309 => x"ffffff",
   6310 => x"ffffff",
   6311 => x"ffffff",
   6312 => x"ffffff",
   6313 => x"ffffff",
   6314 => x"ffffff",
   6315 => x"ffffff",
   6316 => x"ffffff",
   6317 => x"ffffff",
   6318 => x"ffffff",
   6319 => x"ffffff",
   6320 => x"ffffff",
   6321 => x"ffffff",
   6322 => x"ffffff",
   6323 => x"ffffff",
   6324 => x"ffffff",
   6325 => x"ffffff",
   6326 => x"ffffff",
   6327 => x"ffffff",
   6328 => x"ffffff",
   6329 => x"ffffff",
   6330 => x"ffffff",
   6331 => x"ffffff",
   6332 => x"ffffff",
   6333 => x"ffffff",
   6334 => x"ffffff",
   6335 => x"ffffff",
   6336 => x"ffffff",
   6337 => x"ffffff",
   6338 => x"ffffff",
   6339 => x"ffffff",
   6340 => x"ffffff",
   6341 => x"ffffea",
   6342 => x"56afff",
   6343 => x"ffffff",
   6344 => x"ffffff",
   6345 => x"ffffff",
   6346 => x"ffffff",
   6347 => x"ffffff",
   6348 => x"ffffff",
   6349 => x"ffffff",
   6350 => x"ffffff",
   6351 => x"ffffff",
   6352 => x"ffffff",
   6353 => x"ffffff",
   6354 => x"ffffff",
   6355 => x"ffffff",
   6356 => x"ffffff",
   6357 => x"ffffff",
   6358 => x"ffffff",
   6359 => x"ffffff",
   6360 => x"ffffff",
   6361 => x"ffffff",
   6362 => x"ffffff",
   6363 => x"ffffff",
   6364 => x"ffffff",
   6365 => x"ffffff",
   6366 => x"ffffff",
   6367 => x"ffffff",
   6368 => x"ffffff",
   6369 => x"ffffff",
   6370 => x"ffffff",
   6371 => x"ffffff",
   6372 => x"ffffff",
   6373 => x"ffffff",
   6374 => x"ffffff",
   6375 => x"ffffff",
   6376 => x"ffffff",
   6377 => x"ffffff",
   6378 => x"ffffff",
   6379 => x"ffffff",
   6380 => x"ffffff",
   6381 => x"ffffff",
   6382 => x"ffffff",
   6383 => x"ffffff",
   6384 => x"ffffff",
   6385 => x"ffffff",
   6386 => x"ffffff",
   6387 => x"ffffff",
   6388 => x"ffffff",
   6389 => x"ffffff",
   6390 => x"ffffff",
   6391 => x"ffffff",
   6392 => x"ffffff",
   6393 => x"ffffff",
   6394 => x"ffffff",
   6395 => x"ffffff",
   6396 => x"ffffff",
   6397 => x"ffffff",
   6398 => x"ffffff",
   6399 => x"ffffff",
   6400 => x"ffffff",
   6401 => x"ffffff",
   6402 => x"ffffff",
   6403 => x"ffffff",
   6404 => x"ffffff",
   6405 => x"ffffff",
   6406 => x"fffff5",
   6407 => x"c30c30",
   6408 => x"c30c30",
   6409 => x"c30c30",
   6410 => x"c30c30",
   6411 => x"c30c30",
   6412 => x"c30c30",
   6413 => x"c30c30",
   6414 => x"c30c30",
   6415 => x"c30c30",
   6416 => x"c30c30",
   6417 => x"c30c30",
   6418 => x"c30c30",
   6419 => x"c30c30",
   6420 => x"c30c30",
   6421 => x"c30c30",
   6422 => x"c30c30",
   6423 => x"c30c30",
   6424 => x"c30c30",
   6425 => x"c30c30",
   6426 => x"c30c30",
   6427 => x"c30c30",
   6428 => x"c30a2c",
   6429 => x"f3cf3c",
   6430 => x"f3cf3c",
   6431 => x"f3cf3c",
   6432 => x"f3cf3c",
   6433 => x"f3cf3c",
   6434 => x"f3cf3c",
   6435 => x"f3cf3c",
   6436 => x"f3cf3c",
   6437 => x"f3cf3c",
   6438 => x"f3cf3c",
   6439 => x"f3cf1c",
   6440 => x"30c30c",
   6441 => x"30c30c",
   6442 => x"30c30c",
   6443 => x"30c30c",
   6444 => x"30c30c",
   6445 => x"30c30c",
   6446 => x"30c30c",
   6447 => x"30c30c",
   6448 => x"30c30c",
   6449 => x"30c30c",
   6450 => x"30c30c",
   6451 => x"30c30c",
   6452 => x"30c30c",
   6453 => x"30c30c",
   6454 => x"30c30c",
   6455 => x"30c30c",
   6456 => x"30c30c",
   6457 => x"30c30c",
   6458 => x"30c30c",
   6459 => x"30c30c",
   6460 => x"30c30c",
   6461 => x"30c32e",
   6462 => x"ffffff",
   6463 => x"ffffff",
   6464 => x"ffffff",
   6465 => x"ffffff",
   6466 => x"ffffff",
   6467 => x"ffffff",
   6468 => x"ffffff",
   6469 => x"ffffff",
   6470 => x"ffffff",
   6471 => x"ffffff",
   6472 => x"ffffff",
   6473 => x"ffffff",
   6474 => x"ffffff",
   6475 => x"ffffff",
   6476 => x"ffffff",
   6477 => x"ffffff",
   6478 => x"ffffff",
   6479 => x"ffffff",
   6480 => x"ffffff",
   6481 => x"ffffff",
   6482 => x"ffffff",
   6483 => x"ffffff",
   6484 => x"ffffff",
   6485 => x"ffffff",
   6486 => x"ffffff",
   6487 => x"ffffff",
   6488 => x"ffffff",
   6489 => x"ffffff",
   6490 => x"ffffff",
   6491 => x"ffffff",
   6492 => x"ffffff",
   6493 => x"ffffff",
   6494 => x"ffffff",
   6495 => x"ffffff",
   6496 => x"ffffff",
   6497 => x"ffffff",
   6498 => x"ffffff",
   6499 => x"ffffff",
   6500 => x"ffffff",
   6501 => x"fffa95",
   6502 => x"abffff",
   6503 => x"ffffff",
   6504 => x"ffffff",
   6505 => x"ffffff",
   6506 => x"ffffff",
   6507 => x"ffffff",
   6508 => x"ffffff",
   6509 => x"ffffff",
   6510 => x"ffffff",
   6511 => x"ffffff",
   6512 => x"ffffff",
   6513 => x"ffffff",
   6514 => x"ffffff",
   6515 => x"ffffff",
   6516 => x"ffffff",
   6517 => x"ffffff",
   6518 => x"ffffff",
   6519 => x"ffffff",
   6520 => x"ffffff",
   6521 => x"ffffff",
   6522 => x"ffffff",
   6523 => x"ffffff",
   6524 => x"ffffff",
   6525 => x"ffffff",
   6526 => x"ffffff",
   6527 => x"ffffff",
   6528 => x"ffffff",
   6529 => x"ffffff",
   6530 => x"ffffff",
   6531 => x"ffffff",
   6532 => x"ffffff",
   6533 => x"ffffff",
   6534 => x"ffffff",
   6535 => x"ffffff",
   6536 => x"ffffff",
   6537 => x"ffffff",
   6538 => x"ffffff",
   6539 => x"ffffff",
   6540 => x"ffffff",
   6541 => x"ffffff",
   6542 => x"ffffff",
   6543 => x"ffffff",
   6544 => x"ffffff",
   6545 => x"ffffff",
   6546 => x"ffffff",
   6547 => x"ffffff",
   6548 => x"ffffff",
   6549 => x"ffffff",
   6550 => x"ffffff",
   6551 => x"ffffff",
   6552 => x"ffffff",
   6553 => x"ffffff",
   6554 => x"ffffff",
   6555 => x"ffffff",
   6556 => x"ffffff",
   6557 => x"ffffff",
   6558 => x"ffffff",
   6559 => x"ffffff",
   6560 => x"ffffff",
   6561 => x"ffffff",
   6562 => x"ffffff",
   6563 => x"ffffff",
   6564 => x"ffffff",
   6565 => x"ffffff",
   6566 => x"fffd70",
   6567 => x"c30c30",
   6568 => x"c30c30",
   6569 => x"c30c30",
   6570 => x"c30c30",
   6571 => x"c30c30",
   6572 => x"c30c30",
   6573 => x"c30c30",
   6574 => x"c30c30",
   6575 => x"c30c30",
   6576 => x"c30c30",
   6577 => x"c30c30",
   6578 => x"c30c30",
   6579 => x"c30c30",
   6580 => x"c30c30",
   6581 => x"c30c30",
   6582 => x"c30c30",
   6583 => x"c30c30",
   6584 => x"c30c30",
   6585 => x"c30c30",
   6586 => x"c30c30",
   6587 => x"c30c30",
   6588 => x"c28b3c",
   6589 => x"f3cf3c",
   6590 => x"f3cf3c",
   6591 => x"f3cf3c",
   6592 => x"f3cf3c",
   6593 => x"f3cf3c",
   6594 => x"f3cf3c",
   6595 => x"f3cf3c",
   6596 => x"f3cf3c",
   6597 => x"f3cf3c",
   6598 => x"f3cf3c",
   6599 => x"f3cf3c",
   6600 => x"70c30c",
   6601 => x"30c30c",
   6602 => x"30c30c",
   6603 => x"30c30c",
   6604 => x"30c30c",
   6605 => x"30c30c",
   6606 => x"30c30c",
   6607 => x"30c30c",
   6608 => x"30c30c",
   6609 => x"30c30c",
   6610 => x"30c30c",
   6611 => x"30c30c",
   6612 => x"30c30c",
   6613 => x"30c30c",
   6614 => x"30c30c",
   6615 => x"30c30c",
   6616 => x"30c30c",
   6617 => x"30c30c",
   6618 => x"30c30c",
   6619 => x"30c30c",
   6620 => x"30c30c",
   6621 => x"30c30c",
   6622 => x"bbffff",
   6623 => x"ffffff",
   6624 => x"ffffff",
   6625 => x"ffffff",
   6626 => x"ffffff",
   6627 => x"ffffff",
   6628 => x"ffffff",
   6629 => x"ffffff",
   6630 => x"ffffff",
   6631 => x"ffffff",
   6632 => x"ffffff",
   6633 => x"ffffff",
   6634 => x"ffffff",
   6635 => x"ffffff",
   6636 => x"ffffff",
   6637 => x"ffffff",
   6638 => x"ffffff",
   6639 => x"ffffff",
   6640 => x"ffffff",
   6641 => x"ffffff",
   6642 => x"ffffff",
   6643 => x"ffffff",
   6644 => x"ffffff",
   6645 => x"ffffff",
   6646 => x"ffffff",
   6647 => x"ffffff",
   6648 => x"ffffff",
   6649 => x"ffffff",
   6650 => x"ffffff",
   6651 => x"ffffff",
   6652 => x"ffffff",
   6653 => x"ffffff",
   6654 => x"ffffff",
   6655 => x"ffffff",
   6656 => x"ffffff",
   6657 => x"ffffff",
   6658 => x"ffffff",
   6659 => x"ffffff",
   6660 => x"ffffff",
   6661 => x"fea56a",
   6662 => x"ffffff",
   6663 => x"ffffff",
   6664 => x"ffffff",
   6665 => x"ffffff",
   6666 => x"ffffff",
   6667 => x"ffffff",
   6668 => x"ffffff",
   6669 => x"ffffff",
   6670 => x"ffffff",
   6671 => x"ffffff",
   6672 => x"ffffff",
   6673 => x"ffffff",
   6674 => x"ffffff",
   6675 => x"ffffff",
   6676 => x"ffffff",
   6677 => x"ffffff",
   6678 => x"ffffff",
   6679 => x"ffffff",
   6680 => x"ffffff",
   6681 => x"ffffff",
   6682 => x"ffffff",
   6683 => x"ffffff",
   6684 => x"ffffff",
   6685 => x"ffffff",
   6686 => x"ffffff",
   6687 => x"ffffff",
   6688 => x"ffffff",
   6689 => x"ffffff",
   6690 => x"ffffff",
   6691 => x"ffffff",
   6692 => x"ffffff",
   6693 => x"ffffff",
   6694 => x"ffffff",
   6695 => x"ffffff",
   6696 => x"ffffff",
   6697 => x"ffffff",
   6698 => x"ffffff",
   6699 => x"ffffff",
   6700 => x"ffffff",
   6701 => x"ffffff",
   6702 => x"ffffff",
   6703 => x"ffffff",
   6704 => x"ffffff",
   6705 => x"ffffff",
   6706 => x"ffffff",
   6707 => x"ffffff",
   6708 => x"ffffff",
   6709 => x"ffffff",
   6710 => x"ffffff",
   6711 => x"ffffff",
   6712 => x"ffffff",
   6713 => x"ffffff",
   6714 => x"ffffff",
   6715 => x"ffffff",
   6716 => x"ffffff",
   6717 => x"ffffff",
   6718 => x"ffffff",
   6719 => x"ffffff",
   6720 => x"ffffff",
   6721 => x"ffffff",
   6722 => x"ffffff",
   6723 => x"ffffff",
   6724 => x"ffffff",
   6725 => x"ffffff",
   6726 => x"ff5c30",
   6727 => x"c30c30",
   6728 => x"c30c30",
   6729 => x"c30c30",
   6730 => x"c30c30",
   6731 => x"c30c30",
   6732 => x"c30c30",
   6733 => x"c30c30",
   6734 => x"c30c30",
   6735 => x"c30c30",
   6736 => x"c30c30",
   6737 => x"c30c30",
   6738 => x"c30c30",
   6739 => x"c30c30",
   6740 => x"c30c30",
   6741 => x"c30c30",
   6742 => x"c30c30",
   6743 => x"c30c30",
   6744 => x"c30c30",
   6745 => x"c30c30",
   6746 => x"c30c30",
   6747 => x"c30c30",
   6748 => x"92cf3c",
   6749 => x"f3cf3c",
   6750 => x"f3cf3c",
   6751 => x"f3cf3c",
   6752 => x"f3cf3c",
   6753 => x"f3cf3c",
   6754 => x"f3cf3c",
   6755 => x"f3cf3c",
   6756 => x"f3cf3c",
   6757 => x"f3cf3c",
   6758 => x"f3cf3c",
   6759 => x"f3cf3c",
   6760 => x"f1c30c",
   6761 => x"30c30c",
   6762 => x"30c30c",
   6763 => x"30c30c",
   6764 => x"30c30c",
   6765 => x"30c30c",
   6766 => x"30c30c",
   6767 => x"30c30c",
   6768 => x"30c30c",
   6769 => x"30c30c",
   6770 => x"30c30c",
   6771 => x"30c30c",
   6772 => x"30c30c",
   6773 => x"30c30c",
   6774 => x"30c30c",
   6775 => x"30c30c",
   6776 => x"30c30c",
   6777 => x"30c30c",
   6778 => x"30c30c",
   6779 => x"30c30c",
   6780 => x"30c30c",
   6781 => x"30c30c",
   6782 => x"32efff",
   6783 => x"ffffff",
   6784 => x"ffffff",
   6785 => x"ffffff",
   6786 => x"ffffff",
   6787 => x"ffffff",
   6788 => x"ffffff",
   6789 => x"ffffff",
   6790 => x"ffffff",
   6791 => x"ffffff",
   6792 => x"ffffff",
   6793 => x"ffffff",
   6794 => x"ffffff",
   6795 => x"ffffff",
   6796 => x"ffffff",
   6797 => x"ffffff",
   6798 => x"ffffff",
   6799 => x"ffffff",
   6800 => x"ffffff",
   6801 => x"ffffff",
   6802 => x"ffffff",
   6803 => x"ffffff",
   6804 => x"ffffff",
   6805 => x"ffffff",
   6806 => x"ffffff",
   6807 => x"ffffff",
   6808 => x"ffffff",
   6809 => x"ffffff",
   6810 => x"ffffff",
   6811 => x"ffffff",
   6812 => x"ffffff",
   6813 => x"ffffff",
   6814 => x"ffffff",
   6815 => x"ffffff",
   6816 => x"ffffff",
   6817 => x"ffffff",
   6818 => x"ffffff",
   6819 => x"ffffff",
   6820 => x"ffffff",
   6821 => x"a95abf",
   6822 => x"ffffff",
   6823 => x"ffffff",
   6824 => x"ffffff",
   6825 => x"ffffff",
   6826 => x"ffffff",
   6827 => x"ffffff",
   6828 => x"ffffff",
   6829 => x"ffffff",
   6830 => x"ffffff",
   6831 => x"ffffff",
   6832 => x"ffffff",
   6833 => x"ffffff",
   6834 => x"ffffff",
   6835 => x"ffffff",
   6836 => x"ffffff",
   6837 => x"ffffff",
   6838 => x"ffffff",
   6839 => x"ffffff",
   6840 => x"ffffff",
   6841 => x"ffffff",
   6842 => x"ffffff",
   6843 => x"ffffff",
   6844 => x"ffffff",
   6845 => x"ffffff",
   6846 => x"ffffff",
   6847 => x"ffffff",
   6848 => x"ffffff",
   6849 => x"ffffff",
   6850 => x"ffffff",
   6851 => x"ffffff",
   6852 => x"ffffff",
   6853 => x"ffffff",
   6854 => x"ffffff",
   6855 => x"ffffff",
   6856 => x"ffffff",
   6857 => x"ffffff",
   6858 => x"ffffff",
   6859 => x"ffffff",
   6860 => x"ffffff",
   6861 => x"ffffff",
   6862 => x"ffffff",
   6863 => x"ffffff",
   6864 => x"ffffff",
   6865 => x"ffffff",
   6866 => x"ffffff",
   6867 => x"ffffff",
   6868 => x"ffffff",
   6869 => x"ffffff",
   6870 => x"ffffff",
   6871 => x"ffffff",
   6872 => x"ffffff",
   6873 => x"ffffff",
   6874 => x"ffffff",
   6875 => x"ffffff",
   6876 => x"ffffff",
   6877 => x"ffffff",
   6878 => x"ffffff",
   6879 => x"ffffff",
   6880 => x"ffffff",
   6881 => x"ffffff",
   6882 => x"ffffff",
   6883 => x"ffffff",
   6884 => x"ffffff",
   6885 => x"ffffff",
   6886 => x"eb0c30",
   6887 => x"c30c30",
   6888 => x"c30c30",
   6889 => x"c30c30",
   6890 => x"c30c30",
   6891 => x"c30c30",
   6892 => x"c30c30",
   6893 => x"c30c30",
   6894 => x"c30c30",
   6895 => x"c30c30",
   6896 => x"c30c30",
   6897 => x"c30c30",
   6898 => x"c30c30",
   6899 => x"c30c30",
   6900 => x"c30c30",
   6901 => x"c30c30",
   6902 => x"c30c30",
   6903 => x"c30c30",
   6904 => x"c30c30",
   6905 => x"c30c30",
   6906 => x"c30c30",
   6907 => x"c30c24",
   6908 => x"b3cf3c",
   6909 => x"f3cf3c",
   6910 => x"f3cf3c",
   6911 => x"f3cf3c",
   6912 => x"f3cf3c",
   6913 => x"f3cf3c",
   6914 => x"f3cf3c",
   6915 => x"f3cf3c",
   6916 => x"f3cf3c",
   6917 => x"f3cf3c",
   6918 => x"f3cf3c",
   6919 => x"f3cf3c",
   6920 => x"f2c70c",
   6921 => x"30c30c",
   6922 => x"30c30c",
   6923 => x"30c30c",
   6924 => x"30c30c",
   6925 => x"30c30c",
   6926 => x"30c30c",
   6927 => x"30c30c",
   6928 => x"30c30c",
   6929 => x"30c30c",
   6930 => x"30c30c",
   6931 => x"30c30c",
   6932 => x"30c30c",
   6933 => x"30c30c",
   6934 => x"30c30c",
   6935 => x"30c30c",
   6936 => x"30c30c",
   6937 => x"30c30c",
   6938 => x"30c30c",
   6939 => x"30c30c",
   6940 => x"30c30c",
   6941 => x"30c30c",
   6942 => x"31dbbf",
   6943 => x"ffffff",
   6944 => x"ffffff",
   6945 => x"ffffff",
   6946 => x"ffffff",
   6947 => x"ffffff",
   6948 => x"ffffff",
   6949 => x"ffffff",
   6950 => x"ffffff",
   6951 => x"ffffff",
   6952 => x"ffffff",
   6953 => x"ffffff",
   6954 => x"ffffff",
   6955 => x"ffffff",
   6956 => x"ffffff",
   6957 => x"ffffff",
   6958 => x"ffffff",
   6959 => x"ffffff",
   6960 => x"ffffff",
   6961 => x"ffffff",
   6962 => x"ffffff",
   6963 => x"ffffff",
   6964 => x"ffffff",
   6965 => x"ffffff",
   6966 => x"ffffff",
   6967 => x"ffffff",
   6968 => x"ffffff",
   6969 => x"ffffff",
   6970 => x"ffffff",
   6971 => x"ffffff",
   6972 => x"ffffff",
   6973 => x"ffffff",
   6974 => x"ffffff",
   6975 => x"ffffff",
   6976 => x"ffffff",
   6977 => x"ffffff",
   6978 => x"ffffff",
   6979 => x"ffffff",
   6980 => x"ffffea",
   6981 => x"56afff",
   6982 => x"ffffff",
   6983 => x"ffffff",
   6984 => x"ffffff",
   6985 => x"ffffff",
   6986 => x"ffffff",
   6987 => x"ffffff",
   6988 => x"ffffff",
   6989 => x"ffffff",
   6990 => x"ffffff",
   6991 => x"ffffff",
   6992 => x"ffffff",
   6993 => x"ffffff",
   6994 => x"ffffff",
   6995 => x"ffffff",
   6996 => x"ffffff",
   6997 => x"ffffff",
   6998 => x"ffffff",
   6999 => x"ffffff",
   7000 => x"ffffff",
   7001 => x"ffffff",
   7002 => x"ffffff",
   7003 => x"ffffff",
   7004 => x"ffffff",
   7005 => x"ffffff",
   7006 => x"ffffff",
   7007 => x"ffffff",
   7008 => x"ffffff",
   7009 => x"ffffff",
   7010 => x"ffffff",
   7011 => x"ffffff",
   7012 => x"ffffff",
   7013 => x"ffffff",
   7014 => x"ffffff",
   7015 => x"ffffff",
   7016 => x"ffffff",
   7017 => x"ffffff",
   7018 => x"ffffff",
   7019 => x"ffffff",
   7020 => x"ffffff",
   7021 => x"ffffff",
   7022 => x"ffffff",
   7023 => x"ffffff",
   7024 => x"ffffff",
   7025 => x"ffffff",
   7026 => x"ffffff",
   7027 => x"ffffff",
   7028 => x"ffffff",
   7029 => x"ffffff",
   7030 => x"ffffff",
   7031 => x"ffffff",
   7032 => x"ffffff",
   7033 => x"ffffff",
   7034 => x"ffffff",
   7035 => x"ffffff",
   7036 => x"ffffff",
   7037 => x"ffffff",
   7038 => x"ffffff",
   7039 => x"ffffff",
   7040 => x"ffffff",
   7041 => x"ffffff",
   7042 => x"ffffff",
   7043 => x"ffffff",
   7044 => x"ffffff",
   7045 => x"fffffa",
   7046 => x"c30c30",
   7047 => x"c30c30",
   7048 => x"c30c30",
   7049 => x"c30c30",
   7050 => x"c30c30",
   7051 => x"c30c30",
   7052 => x"c30c30",
   7053 => x"c30c30",
   7054 => x"c30c30",
   7055 => x"c30c30",
   7056 => x"c30c30",
   7057 => x"c30c30",
   7058 => x"c30c30",
   7059 => x"c30c30",
   7060 => x"c30c30",
   7061 => x"c30c30",
   7062 => x"c30c30",
   7063 => x"c30c30",
   7064 => x"c30c30",
   7065 => x"c30c30",
   7066 => x"c30c30",
   7067 => x"c3092c",
   7068 => x"f3cf3c",
   7069 => x"f3cf3c",
   7070 => x"f3cf3c",
   7071 => x"f3cf3c",
   7072 => x"f3cf3c",
   7073 => x"f3cf3c",
   7074 => x"f3cf3c",
   7075 => x"f3cf3c",
   7076 => x"f3cf3c",
   7077 => x"f3cf3c",
   7078 => x"f3cf3c",
   7079 => x"f3cf3c",
   7080 => x"f3cb1c",
   7081 => x"30c30c",
   7082 => x"30c30c",
   7083 => x"30c30c",
   7084 => x"30c30c",
   7085 => x"30c30c",
   7086 => x"30c30c",
   7087 => x"30c30c",
   7088 => x"30c30c",
   7089 => x"30c30c",
   7090 => x"30c30c",
   7091 => x"30c30c",
   7092 => x"30c30c",
   7093 => x"30c30c",
   7094 => x"30c30c",
   7095 => x"30c30c",
   7096 => x"30c30c",
   7097 => x"30c30c",
   7098 => x"30c30c",
   7099 => x"30c30c",
   7100 => x"30c30c",
   7101 => x"30c30c",
   7102 => x"30c76e",
   7103 => x"ffffff",
   7104 => x"ffffff",
   7105 => x"ffffff",
   7106 => x"ffffff",
   7107 => x"ffffff",
   7108 => x"ffffff",
   7109 => x"ffffff",
   7110 => x"ffffff",
   7111 => x"ffffff",
   7112 => x"ffffff",
   7113 => x"ffffff",
   7114 => x"ffffff",
   7115 => x"ffffff",
   7116 => x"ffffff",
   7117 => x"ffffff",
   7118 => x"ffffff",
   7119 => x"ffffff",
   7120 => x"ffffff",
   7121 => x"ffffff",
   7122 => x"ffffff",
   7123 => x"ffffff",
   7124 => x"ffffff",
   7125 => x"ffffff",
   7126 => x"ffffff",
   7127 => x"ffffff",
   7128 => x"ffffff",
   7129 => x"ffffff",
   7130 => x"ffffff",
   7131 => x"ffffff",
   7132 => x"ffffff",
   7133 => x"ffffff",
   7134 => x"ffffff",
   7135 => x"ffffff",
   7136 => x"ffffff",
   7137 => x"ffffff",
   7138 => x"ffffff",
   7139 => x"ffffff",
   7140 => x"fffa95",
   7141 => x"abffff",
   7142 => x"ffffff",
   7143 => x"ffffff",
   7144 => x"ffffff",
   7145 => x"ffffff",
   7146 => x"ffffff",
   7147 => x"ffffff",
   7148 => x"ffffff",
   7149 => x"ffffff",
   7150 => x"ffffff",
   7151 => x"ffffff",
   7152 => x"ffffff",
   7153 => x"ffffff",
   7154 => x"ffffff",
   7155 => x"ffffff",
   7156 => x"ffffff",
   7157 => x"ffffff",
   7158 => x"ffffff",
   7159 => x"ffffff",
   7160 => x"ffffff",
   7161 => x"ffffff",
   7162 => x"ffffff",
   7163 => x"ffffff",
   7164 => x"ffffff",
   7165 => x"ffffff",
   7166 => x"ffffff",
   7167 => x"ffffff",
   7168 => x"ffffff",
   7169 => x"ffffff",
   7170 => x"ffffff",
   7171 => x"ffffff",
   7172 => x"ffffff",
   7173 => x"ffffff",
   7174 => x"ffffff",
   7175 => x"ffffff",
   7176 => x"ffffff",
   7177 => x"ffffff",
   7178 => x"ffffff",
   7179 => x"ffffff",
   7180 => x"ffffff",
   7181 => x"ffffff",
   7182 => x"ffffff",
   7183 => x"ffffff",
   7184 => x"ffffff",
   7185 => x"ffffff",
   7186 => x"ffffff",
   7187 => x"ffffff",
   7188 => x"ffffff",
   7189 => x"ffffff",
   7190 => x"ffffff",
   7191 => x"ffffff",
   7192 => x"ffffff",
   7193 => x"ffffff",
   7194 => x"ffffff",
   7195 => x"ffffff",
   7196 => x"ffffff",
   7197 => x"ffffff",
   7198 => x"ffffff",
   7199 => x"ffffff",
   7200 => x"ffffff",
   7201 => x"ffffff",
   7202 => x"ffffff",
   7203 => x"ffffff",
   7204 => x"ffffff",
   7205 => x"fffeb0",
   7206 => x"c30c30",
   7207 => x"c30c30",
   7208 => x"c30c30",
   7209 => x"c30c30",
   7210 => x"c30c30",
   7211 => x"c30c30",
   7212 => x"c30c30",
   7213 => x"c30c30",
   7214 => x"c30c30",
   7215 => x"c30c30",
   7216 => x"c30c30",
   7217 => x"c30c30",
   7218 => x"c30c30",
   7219 => x"c30c30",
   7220 => x"c30c30",
   7221 => x"c30c30",
   7222 => x"c30c30",
   7223 => x"c30c30",
   7224 => x"c30c30",
   7225 => x"c30c30",
   7226 => x"c30c30",
   7227 => x"c24b3c",
   7228 => x"f3cf3c",
   7229 => x"f3cf3c",
   7230 => x"f3cf3c",
   7231 => x"f3cf3c",
   7232 => x"f3cf3c",
   7233 => x"f3cf3c",
   7234 => x"f3cf3c",
   7235 => x"f3cf3c",
   7236 => x"f3cf3c",
   7237 => x"f3cf3c",
   7238 => x"f3cf3c",
   7239 => x"f3cf3c",
   7240 => x"f3cf2c",
   7241 => x"70c30c",
   7242 => x"30c30c",
   7243 => x"30c30c",
   7244 => x"30c30c",
   7245 => x"30c30c",
   7246 => x"30c30c",
   7247 => x"30c30c",
   7248 => x"30c30c",
   7249 => x"30c30c",
   7250 => x"30c30c",
   7251 => x"30c30c",
   7252 => x"30c30c",
   7253 => x"30c30c",
   7254 => x"30c30c",
   7255 => x"30c30c",
   7256 => x"30c30c",
   7257 => x"30c30c",
   7258 => x"30c30c",
   7259 => x"30c30c",
   7260 => x"30c30c",
   7261 => x"30c30c",
   7262 => x"30c31d",
   7263 => x"bbffff",
   7264 => x"ffffff",
   7265 => x"ffffff",
   7266 => x"ffffff",
   7267 => x"ffffff",
   7268 => x"ffffff",
   7269 => x"ffffff",
   7270 => x"ffffff",
   7271 => x"ffffff",
   7272 => x"ffffff",
   7273 => x"ffffff",
   7274 => x"ffffff",
   7275 => x"ffffff",
   7276 => x"ffffff",
   7277 => x"ffffff",
   7278 => x"ffffff",
   7279 => x"ffffff",
   7280 => x"ffffff",
   7281 => x"ffffff",
   7282 => x"ffffff",
   7283 => x"ffffff",
   7284 => x"ffffff",
   7285 => x"ffffff",
   7286 => x"ffffff",
   7287 => x"ffffff",
   7288 => x"ffffff",
   7289 => x"ffffff",
   7290 => x"ffffff",
   7291 => x"ffffff",
   7292 => x"ffffff",
   7293 => x"ffffff",
   7294 => x"ffffff",
   7295 => x"ffffff",
   7296 => x"ffffff",
   7297 => x"ffffff",
   7298 => x"ffffff",
   7299 => x"ffffff",
   7300 => x"fea56a",
   7301 => x"ffffff",
   7302 => x"ffffff",
   7303 => x"ffffff",
   7304 => x"ffffff",
   7305 => x"ffffff",
   7306 => x"ffffff",
   7307 => x"ffffff",
   7308 => x"ffffff",
   7309 => x"ffffff",
   7310 => x"ffffff",
   7311 => x"ffffff",
   7312 => x"ffffff",
   7313 => x"ffffff",
   7314 => x"ffffff",
   7315 => x"ffffff",
   7316 => x"ffffff",
   7317 => x"ffffff",
   7318 => x"ffffff",
   7319 => x"ffffff",
   7320 => x"ffffff",
   7321 => x"ffffff",
   7322 => x"ffffff",
   7323 => x"ffffff",
   7324 => x"ffffff",
   7325 => x"ffffff",
   7326 => x"ffffff",
   7327 => x"ffffff",
   7328 => x"ffffff",
   7329 => x"ffffff",
   7330 => x"ffffff",
   7331 => x"ffffff",
   7332 => x"ffffff",
   7333 => x"ffffff",
   7334 => x"ffffff",
   7335 => x"ffffff",
   7336 => x"ffffff",
   7337 => x"ffffff",
   7338 => x"ffffff",
   7339 => x"ffffff",
   7340 => x"ffffff",
   7341 => x"ffffff",
   7342 => x"ffffff",
   7343 => x"ffffff",
   7344 => x"ffffff",
   7345 => x"ffffff",
   7346 => x"ffffff",
   7347 => x"ffffff",
   7348 => x"ffffff",
   7349 => x"ffffff",
   7350 => x"ffffff",
   7351 => x"ffffff",
   7352 => x"ffffff",
   7353 => x"ffffff",
   7354 => x"ffffff",
   7355 => x"ffffff",
   7356 => x"ffffff",
   7357 => x"ffffff",
   7358 => x"ffffff",
   7359 => x"ffffff",
   7360 => x"ffffff",
   7361 => x"ffffff",
   7362 => x"ffffff",
   7363 => x"ffffff",
   7364 => x"ffffff",
   7365 => x"ffac30",
   7366 => x"c30c30",
   7367 => x"c30c30",
   7368 => x"c30c30",
   7369 => x"c30c30",
   7370 => x"c30c30",
   7371 => x"c30c30",
   7372 => x"c30c30",
   7373 => x"c30c30",
   7374 => x"c30c30",
   7375 => x"c30c30",
   7376 => x"c30c30",
   7377 => x"c30c30",
   7378 => x"c30c30",
   7379 => x"c30c30",
   7380 => x"c30c30",
   7381 => x"c30c30",
   7382 => x"c30c30",
   7383 => x"c30c30",
   7384 => x"c30c30",
   7385 => x"c30c30",
   7386 => x"c30c30",
   7387 => x"c28f3c",
   7388 => x"f3cf3c",
   7389 => x"f3cf3c",
   7390 => x"f3cf3c",
   7391 => x"f3cf3c",
   7392 => x"f3cf3c",
   7393 => x"f3cf3c",
   7394 => x"f3cf3c",
   7395 => x"f3cf3c",
   7396 => x"f3cf3c",
   7397 => x"f3cf3c",
   7398 => x"f3cf3c",
   7399 => x"f3cf3c",
   7400 => x"f3cf3c",
   7401 => x"b0c30c",
   7402 => x"30c30c",
   7403 => x"30c30c",
   7404 => x"30c30c",
   7405 => x"30c30c",
   7406 => x"30c30c",
   7407 => x"30c30c",
   7408 => x"30c30c",
   7409 => x"30c30c",
   7410 => x"30c30c",
   7411 => x"30c30c",
   7412 => x"30c30c",
   7413 => x"30c30c",
   7414 => x"30c30c",
   7415 => x"30c30c",
   7416 => x"30c30c",
   7417 => x"30c30c",
   7418 => x"30c30c",
   7419 => x"30c30c",
   7420 => x"30c30c",
   7421 => x"30c30c",
   7422 => x"30c30c",
   7423 => x"77ffff",
   7424 => x"ffffff",
   7425 => x"ffffff",
   7426 => x"ffffff",
   7427 => x"ffffff",
   7428 => x"ffffff",
   7429 => x"ffffff",
   7430 => x"ffffff",
   7431 => x"ffffff",
   7432 => x"ffffff",
   7433 => x"ffffff",
   7434 => x"ffffff",
   7435 => x"ffffff",
   7436 => x"ffffff",
   7437 => x"ffffff",
   7438 => x"ffffff",
   7439 => x"ffffff",
   7440 => x"ffffff",
   7441 => x"ffffff",
   7442 => x"ffffff",
   7443 => x"ffffff",
   7444 => x"ffffff",
   7445 => x"ffffff",
   7446 => x"ffffff",
   7447 => x"ffffff",
   7448 => x"ffffff",
   7449 => x"ffffff",
   7450 => x"ffffff",
   7451 => x"ffffff",
   7452 => x"ffffff",
   7453 => x"ffffff",
   7454 => x"ffffff",
   7455 => x"ffffff",
   7456 => x"ffffff",
   7457 => x"ffffff",
   7458 => x"ffffff",
   7459 => x"ffffff",
   7460 => x"a95abf",
   7461 => x"ffffff",
   7462 => x"ffffff",
   7463 => x"ffffff",
   7464 => x"ffffff",
   7465 => x"ffffff",
   7466 => x"ffffff",
   7467 => x"ffffff",
   7468 => x"ffffff",
   7469 => x"ffffff",
   7470 => x"ffffff",
   7471 => x"ffffff",
   7472 => x"ffffff",
   7473 => x"ffffff",
   7474 => x"ffffff",
   7475 => x"ffffff",
   7476 => x"ffffff",
   7477 => x"ffffff",
   7478 => x"ffffff",
   7479 => x"ffffff",
   7480 => x"ffffff",
   7481 => x"ffffff",
   7482 => x"ffffff",
   7483 => x"ffffff",
   7484 => x"ffffff",
   7485 => x"ffffff",
   7486 => x"ffffff",
   7487 => x"ffffff",
   7488 => x"ffffff",
   7489 => x"ffffff",
   7490 => x"ffffff",
   7491 => x"ffffff",
   7492 => x"ffffff",
   7493 => x"ffffff",
   7494 => x"ffffff",
   7495 => x"ffffff",
   7496 => x"ffffff",
   7497 => x"ffffff",
   7498 => x"ffffff",
   7499 => x"ffffff",
   7500 => x"ffffff",
   7501 => x"ffffff",
   7502 => x"ffffff",
   7503 => x"ffffff",
   7504 => x"ffffff",
   7505 => x"ffffff",
   7506 => x"ffffff",
   7507 => x"ffffff",
   7508 => x"ffffff",
   7509 => x"ffffff",
   7510 => x"ffffff",
   7511 => x"ffffff",
   7512 => x"ffffff",
   7513 => x"ffffff",
   7514 => x"ffffff",
   7515 => x"ffffff",
   7516 => x"ffffff",
   7517 => x"ffffff",
   7518 => x"ffffff",
   7519 => x"ffffff",
   7520 => x"ffffff",
   7521 => x"ffffff",
   7522 => x"ffffff",
   7523 => x"ffffff",
   7524 => x"ffffff",
   7525 => x"eb5c30",
   7526 => x"c30c30",
   7527 => x"c30c30",
   7528 => x"c30c30",
   7529 => x"c30c30",
   7530 => x"c30c30",
   7531 => x"c30c30",
   7532 => x"c30c30",
   7533 => x"c30c30",
   7534 => x"c30c30",
   7535 => x"c30c30",
   7536 => x"c30c30",
   7537 => x"c30c30",
   7538 => x"c30c30",
   7539 => x"c30c30",
   7540 => x"c30c30",
   7541 => x"c30c30",
   7542 => x"c30c30",
   7543 => x"c30c30",
   7544 => x"c30c30",
   7545 => x"c30c30",
   7546 => x"c30c30",
   7547 => x"a3cf3c",
   7548 => x"f3cf3c",
   7549 => x"f3cf3c",
   7550 => x"f3cf3c",
   7551 => x"f3cf3c",
   7552 => x"f3cf3c",
   7553 => x"f3cf3c",
   7554 => x"f3cf3c",
   7555 => x"f3cf3c",
   7556 => x"f3cf3c",
   7557 => x"f3cf3c",
   7558 => x"f3cf3c",
   7559 => x"f3cf3c",
   7560 => x"f3cf3c",
   7561 => x"f1c30c",
   7562 => x"30c30c",
   7563 => x"30c30c",
   7564 => x"30c30c",
   7565 => x"30c30c",
   7566 => x"30c30c",
   7567 => x"30c30c",
   7568 => x"30c30c",
   7569 => x"30c30c",
   7570 => x"30c30c",
   7571 => x"30c30c",
   7572 => x"30c30c",
   7573 => x"30c30c",
   7574 => x"30c30c",
   7575 => x"30c30c",
   7576 => x"30c30c",
   7577 => x"30c30c",
   7578 => x"30c30c",
   7579 => x"30c30c",
   7580 => x"30c30c",
   7581 => x"30c30c",
   7582 => x"30c30c",
   7583 => x"31dfff",
   7584 => x"ffffff",
   7585 => x"ffffff",
   7586 => x"ffffff",
   7587 => x"ffffff",
   7588 => x"ffffff",
   7589 => x"ffffff",
   7590 => x"ffffff",
   7591 => x"ffffff",
   7592 => x"ffffff",
   7593 => x"ffffff",
   7594 => x"ffffff",
   7595 => x"ffffff",
   7596 => x"ffffff",
   7597 => x"ffffff",
   7598 => x"ffffff",
   7599 => x"ffffff",
   7600 => x"ffffff",
   7601 => x"ffffff",
   7602 => x"ffffff",
   7603 => x"ffffff",
   7604 => x"ffffff",
   7605 => x"ffffff",
   7606 => x"ffffff",
   7607 => x"ffffff",
   7608 => x"ffffff",
   7609 => x"ffffff",
   7610 => x"ffffff",
   7611 => x"ffffff",
   7612 => x"ffffff",
   7613 => x"ffffff",
   7614 => x"ffffff",
   7615 => x"ffffff",
   7616 => x"ffffff",
   7617 => x"ffffff",
   7618 => x"ffffff",
   7619 => x"ffffea",
   7620 => x"56afff",
   7621 => x"ffffff",
   7622 => x"ffffff",
   7623 => x"ffffff",
   7624 => x"ffffff",
   7625 => x"ffffff",
   7626 => x"ffffff",
   7627 => x"ffffff",
   7628 => x"ffffff",
   7629 => x"ffffff",
   7630 => x"ffffff",
   7631 => x"ffffff",
   7632 => x"ffffff",
   7633 => x"ffffff",
   7634 => x"ffffff",
   7635 => x"ffffff",
   7636 => x"ffffff",
   7637 => x"ffffff",
   7638 => x"ffffff",
   7639 => x"ffffff",
   7640 => x"ffffff",
   7641 => x"ffffff",
   7642 => x"ffffff",
   7643 => x"ffffff",
   7644 => x"ffffff",
   7645 => x"ffffff",
   7646 => x"ffffff",
   7647 => x"ffffff",
   7648 => x"ffffff",
   7649 => x"ffffff",
   7650 => x"ffffff",
   7651 => x"ffffff",
   7652 => x"ffffff",
   7653 => x"ffffff",
   7654 => x"ffffff",
   7655 => x"ffffff",
   7656 => x"ffffff",
   7657 => x"ffffff",
   7658 => x"ffffff",
   7659 => x"ffffff",
   7660 => x"ffffff",
   7661 => x"ffffff",
   7662 => x"ffffff",
   7663 => x"ffffff",
   7664 => x"ffffff",
   7665 => x"ffffff",
   7666 => x"ffffff",
   7667 => x"ffffff",
   7668 => x"ffffff",
   7669 => x"ffffff",
   7670 => x"ffffff",
   7671 => x"ffffff",
   7672 => x"ffffff",
   7673 => x"ffffff",
   7674 => x"ffffff",
   7675 => x"ffffff",
   7676 => x"ffffff",
   7677 => x"ffffff",
   7678 => x"ffffff",
   7679 => x"ffffff",
   7680 => x"ffffff",
   7681 => x"ffffff",
   7682 => x"ffffff",
   7683 => x"ffffff",
   7684 => x"ffffff",
   7685 => x"d70c30",
   7686 => x"c30c30",
   7687 => x"c30c30",
   7688 => x"c30c30",
   7689 => x"c30c30",
   7690 => x"c30c30",
   7691 => x"c30c30",
   7692 => x"c30c30",
   7693 => x"c30c30",
   7694 => x"c30c30",
   7695 => x"c30c30",
   7696 => x"c30c30",
   7697 => x"c30c30",
   7698 => x"c30c30",
   7699 => x"c30c30",
   7700 => x"c30c30",
   7701 => x"c30c30",
   7702 => x"c30c30",
   7703 => x"c30c30",
   7704 => x"c30c30",
   7705 => x"c30c30",
   7706 => x"c30c24",
   7707 => x"b3cf3c",
   7708 => x"f3cf3c",
   7709 => x"f3cf3c",
   7710 => x"f3cf3c",
   7711 => x"f3cf3c",
   7712 => x"f3cf3c",
   7713 => x"f3cf3c",
   7714 => x"f3cf3c",
   7715 => x"f3cf3c",
   7716 => x"f3cf3c",
   7717 => x"f3cf3c",
   7718 => x"f3cf3c",
   7719 => x"f3cf3c",
   7720 => x"f3cf3c",
   7721 => x"f3c70c",
   7722 => x"30c30c",
   7723 => x"30c30c",
   7724 => x"30c30c",
   7725 => x"30c30c",
   7726 => x"30c30c",
   7727 => x"30c30c",
   7728 => x"30c30c",
   7729 => x"30c30c",
   7730 => x"30c30c",
   7731 => x"30c30c",
   7732 => x"30c30c",
   7733 => x"30c30c",
   7734 => x"30c30c",
   7735 => x"30c30c",
   7736 => x"30c30c",
   7737 => x"30c30c",
   7738 => x"30c30c",
   7739 => x"30c30c",
   7740 => x"30c30c",
   7741 => x"30c30c",
   7742 => x"30c30c",
   7743 => x"30cbbf",
   7744 => x"ffffff",
   7745 => x"ffffff",
   7746 => x"ffffff",
   7747 => x"ffffff",
   7748 => x"ffffff",
   7749 => x"ffffff",
   7750 => x"ffffff",
   7751 => x"ffffff",
   7752 => x"ffffff",
   7753 => x"ffffff",
   7754 => x"ffffff",
   7755 => x"ffffff",
   7756 => x"ffffff",
   7757 => x"ffffff",
   7758 => x"ffffff",
   7759 => x"ffffff",
   7760 => x"ffffff",
   7761 => x"ffffff",
   7762 => x"ffffff",
   7763 => x"ffffff",
   7764 => x"ffffff",
   7765 => x"ffffff",
   7766 => x"ffffff",
   7767 => x"ffffff",
   7768 => x"ffffff",
   7769 => x"ffffff",
   7770 => x"ffffff",
   7771 => x"ffffff",
   7772 => x"ffffff",
   7773 => x"ffffff",
   7774 => x"ffffff",
   7775 => x"ffffff",
   7776 => x"ffffff",
   7777 => x"ffffff",
   7778 => x"ffffff",
   7779 => x"fffa95",
   7780 => x"abffff",
   7781 => x"ffffff",
   7782 => x"ffffff",
   7783 => x"ffffff",
   7784 => x"ffffff",
   7785 => x"ffffff",
   7786 => x"ffffff",
   7787 => x"ffffff",
   7788 => x"ffffff",
   7789 => x"ffffff",
   7790 => x"ffffff",
   7791 => x"ffffff",
   7792 => x"ffffff",
   7793 => x"ffffff",
   7794 => x"ffffff",
   7795 => x"ffffff",
   7796 => x"ffffff",
   7797 => x"ffffff",
   7798 => x"ffffff",
   7799 => x"ffffff",
   7800 => x"ffffff",
   7801 => x"ffffff",
   7802 => x"ffffff",
   7803 => x"ffffff",
   7804 => x"ffffff",
   7805 => x"ffffff",
   7806 => x"ffffff",
   7807 => x"ffffff",
   7808 => x"ffffff",
   7809 => x"ffffff",
   7810 => x"ffffff",
   7811 => x"ffffff",
   7812 => x"ffffff",
   7813 => x"ffffff",
   7814 => x"ffffff",
   7815 => x"ffffff",
   7816 => x"ffffff",
   7817 => x"ffffff",
   7818 => x"ffffff",
   7819 => x"ffffff",
   7820 => x"ffffff",
   7821 => x"ffffff",
   7822 => x"ffffff",
   7823 => x"ffffff",
   7824 => x"ffffff",
   7825 => x"ffffff",
   7826 => x"ffffff",
   7827 => x"ffffff",
   7828 => x"ffffff",
   7829 => x"ffffff",
   7830 => x"ffffff",
   7831 => x"ffffff",
   7832 => x"ffffff",
   7833 => x"ffffff",
   7834 => x"ffffff",
   7835 => x"ffffff",
   7836 => x"ffffff",
   7837 => x"ffffff",
   7838 => x"ffffff",
   7839 => x"ffffff",
   7840 => x"ffffff",
   7841 => x"ffffff",
   7842 => x"ffffff",
   7843 => x"ffffff",
   7844 => x"fffffa",
   7845 => x"c30c30",
   7846 => x"c30c30",
   7847 => x"c30c30",
   7848 => x"c30c30",
   7849 => x"c30c30",
   7850 => x"c30c30",
   7851 => x"c30c30",
   7852 => x"c30c30",
   7853 => x"c30c30",
   7854 => x"c30c30",
   7855 => x"c30c30",
   7856 => x"c30c30",
   7857 => x"c30c30",
   7858 => x"c30c30",
   7859 => x"c30c30",
   7860 => x"c30c30",
   7861 => x"c30c30",
   7862 => x"c30c30",
   7863 => x"c30c30",
   7864 => x"c30c30",
   7865 => x"c30c30",
   7866 => x"c3092c",
   7867 => x"f3cf3c",
   7868 => x"f3cf3c",
   7869 => x"f3cf3c",
   7870 => x"f3cf3c",
   7871 => x"f3cf3c",
   7872 => x"f3cf3c",
   7873 => x"f3cf3c",
   7874 => x"f3cf3c",
   7875 => x"f3cf3c",
   7876 => x"f3cf3c",
   7877 => x"f3cf3c",
   7878 => x"f3cf3c",
   7879 => x"f3cf3c",
   7880 => x"f3cf3c",
   7881 => x"f3cb1c",
   7882 => x"30c30c",
   7883 => x"30c30c",
   7884 => x"30c30c",
   7885 => x"30c30c",
   7886 => x"30c30c",
   7887 => x"30c30c",
   7888 => x"30c30c",
   7889 => x"30c30c",
   7890 => x"30c30c",
   7891 => x"30c30c",
   7892 => x"30c30c",
   7893 => x"30c30c",
   7894 => x"30c30c",
   7895 => x"30c30c",
   7896 => x"30c30c",
   7897 => x"30c30c",
   7898 => x"30c30c",
   7899 => x"30c30c",
   7900 => x"30c30c",
   7901 => x"30c30c",
   7902 => x"30c30c",
   7903 => x"30c76e",
   7904 => x"ffffff",
   7905 => x"ffffff",
   7906 => x"ffffff",
   7907 => x"ffffff",
   7908 => x"ffffff",
   7909 => x"ffffff",
   7910 => x"ffffff",
   7911 => x"ffffff",
   7912 => x"ffffff",
   7913 => x"ffffff",
   7914 => x"ffffff",
   7915 => x"ffffff",
   7916 => x"ffffff",
   7917 => x"ffffff",
   7918 => x"ffffff",
   7919 => x"ffffff",
   7920 => x"ffffff",
   7921 => x"ffffff",
   7922 => x"ffffff",
   7923 => x"ffffff",
   7924 => x"ffffff",
   7925 => x"ffffff",
   7926 => x"ffffff",
   7927 => x"ffffff",
   7928 => x"ffffff",
   7929 => x"ffffff",
   7930 => x"ffffff",
   7931 => x"ffffff",
   7932 => x"ffffff",
   7933 => x"ffffff",
   7934 => x"ffffff",
   7935 => x"ffffff",
   7936 => x"ffffff",
   7937 => x"ffffff",
   7938 => x"ffffff",
   7939 => x"fea56a",
   7940 => x"ffffff",
   7941 => x"ffffff",
   7942 => x"ffffff",
   7943 => x"ffffff",
   7944 => x"ffffff",
   7945 => x"ffffff",
   7946 => x"ffffff",
   7947 => x"ffffff",
   7948 => x"ffffff",
   7949 => x"ffffff",
   7950 => x"ffffff",
   7951 => x"ffffff",
   7952 => x"ffffff",
   7953 => x"ffffff",
   7954 => x"ffffff",
   7955 => x"ffffff",
   7956 => x"ffffff",
   7957 => x"ffffff",
   7958 => x"ffffff",
   7959 => x"ffffff",
   7960 => x"ffffff",
   7961 => x"ffffff",
   7962 => x"ffffff",
   7963 => x"ffffff",
   7964 => x"ffffff",
   7965 => x"ffffff",
   7966 => x"ffffff",
   7967 => x"ffffff",
   7968 => x"ffffff",
   7969 => x"ffffff",
   7970 => x"ffffff",
   7971 => x"ffffff",
   7972 => x"ffffff",
   7973 => x"ffffff",
   7974 => x"ffffff",
   7975 => x"ffffff",
   7976 => x"ffffff",
   7977 => x"ffffff",
   7978 => x"ffffff",
   7979 => x"ffffff",
   7980 => x"ffffff",
   7981 => x"ffffff",
   7982 => x"ffffff",
   7983 => x"ffffff",
   7984 => x"ffffff",
   7985 => x"ffffff",
   7986 => x"ffffff",
   7987 => x"ffffff",
   7988 => x"ffffff",
   7989 => x"ffffff",
   7990 => x"ffffff",
   7991 => x"ffffff",
   7992 => x"ffffff",
   7993 => x"ffffff",
   7994 => x"ffffff",
   7995 => x"ffffff",
   7996 => x"ffffff",
   7997 => x"ffffff",
   7998 => x"ffffff",
   7999 => x"ffffff",
   8000 => x"ffffff",
   8001 => x"ffffff",
   8002 => x"ffffff",
   8003 => x"ffffff",
   8004 => x"fffeb0",
   8005 => x"c30c30",
   8006 => x"c30c30",
   8007 => x"c30c30",
   8008 => x"c30c30",
   8009 => x"c30c30",
   8010 => x"c30c30",
   8011 => x"c30c30",
   8012 => x"c30c30",
   8013 => x"c30c30",
   8014 => x"c30c30",
   8015 => x"c30c30",
   8016 => x"c30c30",
   8017 => x"c30c30",
   8018 => x"c30c30",
   8019 => x"c30c30",
   8020 => x"c30c30",
   8021 => x"c30c30",
   8022 => x"c30c30",
   8023 => x"c30c30",
   8024 => x"c30c30",
   8025 => x"c30c30",
   8026 => x"c3063c",
   8027 => x"f3cf3c",
   8028 => x"f3cf3c",
   8029 => x"f3cf3c",
   8030 => x"f3cf3c",
   8031 => x"f3cf3c",
   8032 => x"f3cf3c",
   8033 => x"f3cf3c",
   8034 => x"f3cf3c",
   8035 => x"f3cf3c",
   8036 => x"f3cf3c",
   8037 => x"f3cf3c",
   8038 => x"f3cf3c",
   8039 => x"f3cf3c",
   8040 => x"f3cf3c",
   8041 => x"f3cf2c",
   8042 => x"30c30c",
   8043 => x"30c30c",
   8044 => x"30c30c",
   8045 => x"30c30c",
   8046 => x"30c30c",
   8047 => x"30c30c",
   8048 => x"30c30c",
   8049 => x"30c30c",
   8050 => x"30c30c",
   8051 => x"30c30c",
   8052 => x"30c30c",
   8053 => x"30c30c",
   8054 => x"30c30c",
   8055 => x"30c30c",
   8056 => x"30c30c",
   8057 => x"30c30c",
   8058 => x"30c30c",
   8059 => x"30c30c",
   8060 => x"30c30c",
   8061 => x"30c30c",
   8062 => x"30c30c",
   8063 => x"30c31d",
   8064 => x"ffffff",
   8065 => x"ffffff",
   8066 => x"ffffff",
   8067 => x"ffffff",
   8068 => x"ffffff",
   8069 => x"ffffff",
   8070 => x"ffffff",
   8071 => x"ffffff",
   8072 => x"ffffff",
   8073 => x"ffffff",
   8074 => x"ffffff",
   8075 => x"ffffff",
   8076 => x"ffffff",
   8077 => x"ffffff",
   8078 => x"ffffff",
   8079 => x"ffffff",
   8080 => x"ffffff",
   8081 => x"ffffff",
   8082 => x"ffffff",
   8083 => x"ffffff",
   8084 => x"ffffff",
   8085 => x"ffffff",
   8086 => x"ffffff",
   8087 => x"ffffff",
   8088 => x"ffffff",
   8089 => x"ffffff",
   8090 => x"ffffff",
   8091 => x"ffffff",
   8092 => x"ffffff",
   8093 => x"ffffff",
   8094 => x"ffffff",
   8095 => x"ffffff",
   8096 => x"ffffff",
   8097 => x"ffffff",
   8098 => x"ffffff",
   8099 => x"a95abf",
   8100 => x"ffffff",
   8101 => x"ffffff",
   8102 => x"ffffff",
   8103 => x"ffffff",
   8104 => x"ffffff",
   8105 => x"ffffff",
   8106 => x"ffffff",
   8107 => x"ffffff",
   8108 => x"ffffff",
   8109 => x"ffffff",
   8110 => x"ffffff",
   8111 => x"ffffff",
   8112 => x"ffffff",
   8113 => x"ffffff",
   8114 => x"ffffff",
   8115 => x"ffffff",
   8116 => x"ffffff",
   8117 => x"ffffff",
   8118 => x"ffffff",
   8119 => x"ffffff",
   8120 => x"ffffff",
   8121 => x"ffffff",
   8122 => x"ffffff",
   8123 => x"ffffff",
   8124 => x"ffffff",
   8125 => x"ffffff",
   8126 => x"ffffff",
   8127 => x"ffffff",
   8128 => x"ffffff",
   8129 => x"ffffff",
   8130 => x"ffffff",
   8131 => x"ffffff",
   8132 => x"ffffff",
   8133 => x"ffffff",
   8134 => x"ffffff",
   8135 => x"ffffff",
   8136 => x"ffffff",
   8137 => x"ffffff",
   8138 => x"ffffff",
   8139 => x"ffffff",
   8140 => x"ffffff",
   8141 => x"ffffff",
   8142 => x"ffffff",
   8143 => x"ffffff",
   8144 => x"ffffff",
   8145 => x"ffffff",
   8146 => x"ffffff",
   8147 => x"ffffff",
   8148 => x"ffffff",
   8149 => x"ffffff",
   8150 => x"ffffff",
   8151 => x"ffffff",
   8152 => x"ffffff",
   8153 => x"ffffff",
   8154 => x"ffffff",
   8155 => x"ffffff",
   8156 => x"ffffff",
   8157 => x"ffffff",
   8158 => x"ffffff",
   8159 => x"ffffff",
   8160 => x"ffffff",
   8161 => x"ffffff",
   8162 => x"ffffff",
   8163 => x"ffffff",
   8164 => x"ffad70",
   8165 => x"c30c30",
   8166 => x"c30c30",
   8167 => x"c30c30",
   8168 => x"c30c30",
   8169 => x"c30c30",
   8170 => x"c30c30",
   8171 => x"c30c30",
   8172 => x"c30c30",
   8173 => x"c30c30",
   8174 => x"c30c30",
   8175 => x"c30c30",
   8176 => x"c30c30",
   8177 => x"c30c30",
   8178 => x"c30c30",
   8179 => x"c30c30",
   8180 => x"c30c30",
   8181 => x"c30c30",
   8182 => x"c30c30",
   8183 => x"c30c30",
   8184 => x"c30c30",
   8185 => x"c30c30",
   8186 => x"c28f3c",
   8187 => x"f3cf3c",
   8188 => x"f3cf3c",
   8189 => x"f3cf3c",
   8190 => x"f3cf3c",
   8191 => x"f3cf3c",
   8192 => x"f3cf3c",
   8193 => x"f3cf3c",
   8194 => x"f3cf3c",
   8195 => x"f3cf3c",
   8196 => x"f3cf3c",
   8197 => x"f3cf3c",
   8198 => x"f3cf3c",
   8199 => x"f3cf3c",
   8200 => x"f3cf3c",
   8201 => x"f3cf3c",
   8202 => x"70c30c",
   8203 => x"30c30c",
   8204 => x"30c30c",
   8205 => x"30c30c",
   8206 => x"30c30c",
   8207 => x"30c30c",
   8208 => x"30c30c",
   8209 => x"30c30c",
   8210 => x"30c30c",
   8211 => x"30c30c",
   8212 => x"30c30c",
   8213 => x"30c30c",
   8214 => x"30c30c",
   8215 => x"30c30c",
   8216 => x"30c30c",
   8217 => x"30c30c",
   8218 => x"30c30c",
   8219 => x"30c30c",
   8220 => x"30c30c",
   8221 => x"30c30c",
   8222 => x"30c30c",
   8223 => x"30c30c",
   8224 => x"77ffff",
   8225 => x"ffffff",
   8226 => x"ffffff",
   8227 => x"ffffff",
   8228 => x"ffffff",
   8229 => x"ffffff",
   8230 => x"ffffff",
   8231 => x"ffffff",
   8232 => x"ffffff",
   8233 => x"ffffff",
   8234 => x"ffffff",
   8235 => x"ffffff",
   8236 => x"ffffff",
   8237 => x"ffffff",
   8238 => x"ffffff",
   8239 => x"ffffff",
   8240 => x"ffffff",
   8241 => x"ffffff",
   8242 => x"ffffff",
   8243 => x"ffffff",
   8244 => x"ffffff",
   8245 => x"ffffff",
   8246 => x"ffffff",
   8247 => x"ffffff",
   8248 => x"ffffff",
   8249 => x"ffffff",
   8250 => x"ffffff",
   8251 => x"ffffff",
   8252 => x"ffffff",
   8253 => x"ffffff",
   8254 => x"ffffff",
   8255 => x"ffffff",
   8256 => x"ffffff",
   8257 => x"ffffff",
   8258 => x"ffffea",
   8259 => x"56afff",
   8260 => x"ffffff",
   8261 => x"ffffff",
   8262 => x"ffffff",
   8263 => x"ffffff",
   8264 => x"ffffff",
   8265 => x"ffffff",
   8266 => x"ffffff",
   8267 => x"ffffff",
   8268 => x"ffffff",
   8269 => x"ffffff",
   8270 => x"ffffff",
   8271 => x"ffffff",
   8272 => x"ffffff",
   8273 => x"ffffff",
   8274 => x"ffffff",
   8275 => x"ffffff",
   8276 => x"ffffff",
   8277 => x"ffffff",
   8278 => x"ffffff",
   8279 => x"ffffff",
   8280 => x"ffffff",
   8281 => x"ffffff",
   8282 => x"ffffff",
   8283 => x"ffffff",
   8284 => x"ffffff",
   8285 => x"ffffff",
   8286 => x"ffffff",
   8287 => x"ffffff",
   8288 => x"ffffff",
   8289 => x"ffffff",
   8290 => x"ffffff",
   8291 => x"ffffff",
   8292 => x"ffffff",
   8293 => x"ffffff",
   8294 => x"ffffff",
   8295 => x"ffffff",
   8296 => x"ffffff",
   8297 => x"ffffff",
   8298 => x"ffffff",
   8299 => x"ffffff",
   8300 => x"ffffff",
   8301 => x"ffffff",
   8302 => x"ffffff",
   8303 => x"ffffff",
   8304 => x"ffffff",
   8305 => x"ffffff",
   8306 => x"ffffff",
   8307 => x"ffffff",
   8308 => x"ffffff",
   8309 => x"ffffff",
   8310 => x"ffffff",
   8311 => x"ffffff",
   8312 => x"ffffff",
   8313 => x"ffffff",
   8314 => x"ffffff",
   8315 => x"ffffff",
   8316 => x"ffffff",
   8317 => x"ffffff",
   8318 => x"ffffff",
   8319 => x"ffffff",
   8320 => x"ffffff",
   8321 => x"ffffff",
   8322 => x"ffffff",
   8323 => x"ffffff",
   8324 => x"ff5c30",
   8325 => x"c30c30",
   8326 => x"c30c30",
   8327 => x"c30c30",
   8328 => x"c30c30",
   8329 => x"c30c30",
   8330 => x"c30c30",
   8331 => x"c30c30",
   8332 => x"c30c30",
   8333 => x"c30c30",
   8334 => x"c30c30",
   8335 => x"c30c30",
   8336 => x"c30c30",
   8337 => x"c30c30",
   8338 => x"c30c30",
   8339 => x"c30c30",
   8340 => x"c30c30",
   8341 => x"c30c30",
   8342 => x"c30c30",
   8343 => x"c30c30",
   8344 => x"c30c30",
   8345 => x"c30c30",
   8346 => x"92cf3c",
   8347 => x"f3cf3c",
   8348 => x"f3cf3c",
   8349 => x"f3cf3c",
   8350 => x"f3cf3c",
   8351 => x"f3cf3c",
   8352 => x"f3cf3c",
   8353 => x"f3cf3c",
   8354 => x"f3cf3c",
   8355 => x"f3cf3c",
   8356 => x"f3cf3c",
   8357 => x"f3cf3c",
   8358 => x"f3cf3c",
   8359 => x"f3cf3c",
   8360 => x"f3cf3c",
   8361 => x"f3cf3c",
   8362 => x"f1c30c",
   8363 => x"30c30c",
   8364 => x"30c30c",
   8365 => x"30c30c",
   8366 => x"30c30c",
   8367 => x"30c30c",
   8368 => x"30c30c",
   8369 => x"30c30c",
   8370 => x"30c30c",
   8371 => x"30c30c",
   8372 => x"30c30c",
   8373 => x"30c30c",
   8374 => x"30c30c",
   8375 => x"30c30c",
   8376 => x"30c30c",
   8377 => x"30c30c",
   8378 => x"30c30c",
   8379 => x"30c30c",
   8380 => x"30c30c",
   8381 => x"30c30c",
   8382 => x"30c30c",
   8383 => x"30c30c",
   8384 => x"32efff",
   8385 => x"ffffff",
   8386 => x"ffffff",
   8387 => x"ffffff",
   8388 => x"ffffff",
   8389 => x"ffffff",
   8390 => x"ffffff",
   8391 => x"ffffff",
   8392 => x"ffffff",
   8393 => x"ffffff",
   8394 => x"ffffff",
   8395 => x"ffffff",
   8396 => x"ffffff",
   8397 => x"ffffff",
   8398 => x"ffffff",
   8399 => x"ffffff",
   8400 => x"ffffff",
   8401 => x"ffffff",
   8402 => x"ffffff",
   8403 => x"ffffff",
   8404 => x"ffffff",
   8405 => x"ffffff",
   8406 => x"ffffff",
   8407 => x"ffffff",
   8408 => x"ffffff",
   8409 => x"ffffff",
   8410 => x"ffffff",
   8411 => x"ffffff",
   8412 => x"ffffff",
   8413 => x"ffffff",
   8414 => x"ffffff",
   8415 => x"ffffff",
   8416 => x"ffffff",
   8417 => x"ffffff",
   8418 => x"fffa95",
   8419 => x"abffff",
   8420 => x"ffffff",
   8421 => x"ffffff",
   8422 => x"ffffff",
   8423 => x"ffffff",
   8424 => x"ffffff",
   8425 => x"ffffff",
   8426 => x"ffffff",
   8427 => x"ffffff",
   8428 => x"ffffff",
   8429 => x"ffffff",
   8430 => x"ffffff",
   8431 => x"ffffff",
   8432 => x"ffffff",
   8433 => x"ffffff",
   8434 => x"ffffff",
   8435 => x"ffffff",
   8436 => x"ffffff",
   8437 => x"ffffff",
   8438 => x"ffffff",
   8439 => x"ffffff",
   8440 => x"ffffff",
   8441 => x"ffffff",
   8442 => x"ffffff",
   8443 => x"ffffff",
   8444 => x"ffffff",
   8445 => x"ffffff",
   8446 => x"ffffff",
   8447 => x"ffffff",
   8448 => x"ffffff",
   8449 => x"ffffff",
   8450 => x"ffffff",
   8451 => x"ffffff",
   8452 => x"ffffff",
   8453 => x"ffffff",
   8454 => x"ffffff",
   8455 => x"ffffff",
   8456 => x"ffffff",
   8457 => x"ffffff",
   8458 => x"ffffff",
   8459 => x"ffffff",
   8460 => x"ffffff",
   8461 => x"ffffff",
   8462 => x"ffffff",
   8463 => x"ffffff",
   8464 => x"ffffff",
   8465 => x"ffffff",
   8466 => x"ffffff",
   8467 => x"ffffff",
   8468 => x"ffffff",
   8469 => x"ffffff",
   8470 => x"ffffff",
   8471 => x"ffffff",
   8472 => x"ffffff",
   8473 => x"ffffff",
   8474 => x"ffffff",
   8475 => x"ffffff",
   8476 => x"ffffff",
   8477 => x"ffffff",
   8478 => x"ffffff",
   8479 => x"ffffff",
   8480 => x"ffffff",
   8481 => x"ffffff",
   8482 => x"ffffff",
   8483 => x"ffffff",
   8484 => x"eb0c30",
   8485 => x"c30c30",
   8486 => x"c30c30",
   8487 => x"c30c30",
   8488 => x"c30c30",
   8489 => x"c30c30",
   8490 => x"c30c30",
   8491 => x"c30c30",
   8492 => x"c30c30",
   8493 => x"c30c30",
   8494 => x"c30c30",
   8495 => x"c30c30",
   8496 => x"c30c30",
   8497 => x"c30c30",
   8498 => x"c30c30",
   8499 => x"c30c30",
   8500 => x"c30c30",
   8501 => x"c30c30",
   8502 => x"c30c30",
   8503 => x"c30c30",
   8504 => x"c30c30",
   8505 => x"c30c34",
   8506 => x"73cf3c",
   8507 => x"f3cf3c",
   8508 => x"f3cf3c",
   8509 => x"f3cf3c",
   8510 => x"f3cf3c",
   8511 => x"f3cf3c",
   8512 => x"f3cf3c",
   8513 => x"f3cf3c",
   8514 => x"f3cf3c",
   8515 => x"f3cf3c",
   8516 => x"f3cf3c",
   8517 => x"f3cf3c",
   8518 => x"f3cf3c",
   8519 => x"f3cf3c",
   8520 => x"f3cf3c",
   8521 => x"f3cf3c",
   8522 => x"f2c70c",
   8523 => x"30c30c",
   8524 => x"30c30c",
   8525 => x"30c30c",
   8526 => x"30c30c",
   8527 => x"30c30c",
   8528 => x"30c30c",
   8529 => x"30c30c",
   8530 => x"30c30c",
   8531 => x"30c30c",
   8532 => x"30c30c",
   8533 => x"30c30c",
   8534 => x"30c30c",
   8535 => x"30c30c",
   8536 => x"30c30c",
   8537 => x"30c30c",
   8538 => x"30c30c",
   8539 => x"30c30c",
   8540 => x"30c30c",
   8541 => x"30c30c",
   8542 => x"30c30c",
   8543 => x"30c30c",
   8544 => x"31dbbf",
   8545 => x"ffffff",
   8546 => x"ffffff",
   8547 => x"ffffff",
   8548 => x"ffffff",
   8549 => x"ffffff",
   8550 => x"ffffff",
   8551 => x"ffffff",
   8552 => x"ffffff",
   8553 => x"ffffff",
   8554 => x"ffffff",
   8555 => x"ffffff",
   8556 => x"ffffff",
   8557 => x"ffffff",
   8558 => x"ffffff",
   8559 => x"ffffff",
   8560 => x"ffffff",
   8561 => x"ffffff",
   8562 => x"ffffff",
   8563 => x"ffffff",
   8564 => x"ffffff",
   8565 => x"ffffff",
   8566 => x"ffffff",
   8567 => x"ffffff",
   8568 => x"ffffff",
   8569 => x"ffffff",
   8570 => x"ffffff",
   8571 => x"ffffff",
   8572 => x"ffffff",
   8573 => x"ffffff",
   8574 => x"ffffff",
   8575 => x"ffffff",
   8576 => x"ffffff",
   8577 => x"ffffff",
   8578 => x"fea56a",
   8579 => x"ffffff",
   8580 => x"ffffff",
   8581 => x"ffffff",
   8582 => x"ffffff",
   8583 => x"ffffff",
   8584 => x"ffffff",
   8585 => x"ffffff",
   8586 => x"ffffff",
   8587 => x"ffffff",
   8588 => x"ffffff",
   8589 => x"ffffff",
   8590 => x"ffffff",
   8591 => x"ffffff",
   8592 => x"ffffff",
   8593 => x"ffffff",
   8594 => x"ffffff",
   8595 => x"ffffff",
   8596 => x"ffffff",
   8597 => x"ffffff",
   8598 => x"ffffff",
   8599 => x"ffffff",
   8600 => x"ffffff",
   8601 => x"ffffff",
   8602 => x"ffffff",
   8603 => x"ffffff",
   8604 => x"ffffff",
   8605 => x"ffffff",
   8606 => x"ffffff",
   8607 => x"ffffff",
   8608 => x"ffffff",
   8609 => x"ffffff",
   8610 => x"ffffff",
   8611 => x"ffffff",
   8612 => x"ffffff",
   8613 => x"ffffff",
   8614 => x"ffffff",
   8615 => x"ffffff",
   8616 => x"ffffff",
   8617 => x"ffffff",
   8618 => x"ffffff",
   8619 => x"ffffff",
   8620 => x"ffffff",
   8621 => x"ffffff",
   8622 => x"ffffff",
   8623 => x"ffffff",
   8624 => x"ffffff",
   8625 => x"ffffff",
   8626 => x"ffffff",
   8627 => x"ffffff",
   8628 => x"ffffff",
   8629 => x"ffffff",
   8630 => x"ffffff",
   8631 => x"ffffff",
   8632 => x"ffffff",
   8633 => x"ffffff",
   8634 => x"ffffff",
   8635 => x"ffffff",
   8636 => x"ffffff",
   8637 => x"ffffff",
   8638 => x"ffffff",
   8639 => x"ffffff",
   8640 => x"ffffff",
   8641 => x"ffffff",
   8642 => x"ffffff",
   8643 => x"fffffa",
   8644 => x"d70c30",
   8645 => x"c30c30",
   8646 => x"c30c30",
   8647 => x"c30c30",
   8648 => x"c30c30",
   8649 => x"c30c30",
   8650 => x"c30c30",
   8651 => x"c30c30",
   8652 => x"c30c30",
   8653 => x"c30c30",
   8654 => x"c30c30",
   8655 => x"c30c30",
   8656 => x"c30c30",
   8657 => x"c30c30",
   8658 => x"c30c30",
   8659 => x"c30c30",
   8660 => x"c30c30",
   8661 => x"c30c30",
   8662 => x"c30c30",
   8663 => x"c30c30",
   8664 => x"c30c30",
   8665 => x"c30c28",
   8666 => x"f3cf3c",
   8667 => x"f3cf3c",
   8668 => x"f3cf3c",
   8669 => x"f3cf3c",
   8670 => x"f3cf3c",
   8671 => x"f3cf3c",
   8672 => x"f3cf3c",
   8673 => x"f3cf3c",
   8674 => x"f3cf3c",
   8675 => x"f3cf3c",
   8676 => x"f3cf3c",
   8677 => x"f3cf3c",
   8678 => x"f3cf3c",
   8679 => x"f3cf3c",
   8680 => x"f3cf3c",
   8681 => x"f3cf3c",
   8682 => x"f3c70c",
   8683 => x"30c30c",
   8684 => x"30c30c",
   8685 => x"30c30c",
   8686 => x"30c30c",
   8687 => x"30c30c",
   8688 => x"30c30c",
   8689 => x"30c30c",
   8690 => x"30c30c",
   8691 => x"30c30c",
   8692 => x"30c30c",
   8693 => x"30c30c",
   8694 => x"30c30c",
   8695 => x"30c30c",
   8696 => x"30c30c",
   8697 => x"30c30c",
   8698 => x"30c30c",
   8699 => x"30c30c",
   8700 => x"30c30c",
   8701 => x"30c30c",
   8702 => x"30c30c",
   8703 => x"30c30c",
   8704 => x"30c77f",
   8705 => x"ffffff",
   8706 => x"ffffff",
   8707 => x"ffffff",
   8708 => x"ffffff",
   8709 => x"ffffff",
   8710 => x"ffffff",
   8711 => x"ffffff",
   8712 => x"ffffff",
   8713 => x"ffffff",
   8714 => x"ffffff",
   8715 => x"ffffff",
   8716 => x"ffffff",
   8717 => x"ffffff",
   8718 => x"ffffff",
   8719 => x"ffffff",
   8720 => x"ffffff",
   8721 => x"ffffff",
   8722 => x"ffffff",
   8723 => x"ffffff",
   8724 => x"ffffff",
   8725 => x"ffffff",
   8726 => x"ffffff",
   8727 => x"ffffff",
   8728 => x"ffffff",
   8729 => x"ffffff",
   8730 => x"ffffff",
   8731 => x"ffffff",
   8732 => x"ffffff",
   8733 => x"ffffff",
   8734 => x"ffffff",
   8735 => x"ffffff",
   8736 => x"ffffff",
   8737 => x"ffffff",
   8738 => x"a95abf",
   8739 => x"ffffff",
   8740 => x"ffffff",
   8741 => x"ffffff",
   8742 => x"ffffff",
   8743 => x"ffffff",
   8744 => x"ffffff",
   8745 => x"ffffff",
   8746 => x"ffffff",
   8747 => x"ffffff",
   8748 => x"ffffff",
   8749 => x"ffffff",
   8750 => x"ffffff",
   8751 => x"ffffff",
   8752 => x"ffffff",
   8753 => x"ffffff",
   8754 => x"ffffff",
   8755 => x"ffffff",
   8756 => x"ffffff",
   8757 => x"ffffff",
   8758 => x"ffffff",
   8759 => x"ffffff",
   8760 => x"ffffff",
   8761 => x"ffffff",
   8762 => x"ffffff",
   8763 => x"ffffff",
   8764 => x"ffffff",
   8765 => x"ffffff",
   8766 => x"ffffff",
   8767 => x"ffffff",
   8768 => x"ffffff",
   8769 => x"ffffff",
   8770 => x"ffffff",
   8771 => x"ffffff",
   8772 => x"ffffff",
   8773 => x"ffffff",
   8774 => x"ffffff",
   8775 => x"ffffff",
   8776 => x"ffffff",
   8777 => x"ffffff",
   8778 => x"ffffff",
   8779 => x"ffffff",
   8780 => x"ffffff",
   8781 => x"ffffff",
   8782 => x"ffffff",
   8783 => x"ffffff",
   8784 => x"ffffff",
   8785 => x"ffffff",
   8786 => x"ffffff",
   8787 => x"ffffff",
   8788 => x"ffffff",
   8789 => x"ffffff",
   8790 => x"ffffff",
   8791 => x"ffffff",
   8792 => x"ffffff",
   8793 => x"ffffff",
   8794 => x"ffffff",
   8795 => x"ffffff",
   8796 => x"ffffff",
   8797 => x"ffffff",
   8798 => x"ffffff",
   8799 => x"ffffff",
   8800 => x"ffffff",
   8801 => x"ffffff",
   8802 => x"ffffff",
   8803 => x"fffff5",
   8804 => x"c30c30",
   8805 => x"c30c30",
   8806 => x"c30c30",
   8807 => x"c30c30",
   8808 => x"c30c30",
   8809 => x"c30c30",
   8810 => x"c30c30",
   8811 => x"c30c30",
   8812 => x"c30c30",
   8813 => x"c30c30",
   8814 => x"c30c30",
   8815 => x"c30c30",
   8816 => x"c30c30",
   8817 => x"c30c30",
   8818 => x"c30c30",
   8819 => x"c30c30",
   8820 => x"c30c30",
   8821 => x"c30c30",
   8822 => x"c30c30",
   8823 => x"c30c30",
   8824 => x"c30c30",
   8825 => x"c3092c",
   8826 => x"f3cf3c",
   8827 => x"f3cf3c",
   8828 => x"f3cf3c",
   8829 => x"f3cf3c",
   8830 => x"f3cf3c",
   8831 => x"f3cf3c",
   8832 => x"f3cf3c",
   8833 => x"f3cf3c",
   8834 => x"f3cf3c",
   8835 => x"f3cf3c",
   8836 => x"f3cf3c",
   8837 => x"f3cf3c",
   8838 => x"f3cf3c",
   8839 => x"f3cf3c",
   8840 => x"f3cf3c",
   8841 => x"f3cf3c",
   8842 => x"f3cf1c",
   8843 => x"30c30c",
   8844 => x"30c30c",
   8845 => x"30c30c",
   8846 => x"30c30c",
   8847 => x"30c30c",
   8848 => x"30c30c",
   8849 => x"30c30c",
   8850 => x"30c30c",
   8851 => x"30c30c",
   8852 => x"30c30c",
   8853 => x"30c30c",
   8854 => x"30c30c",
   8855 => x"30c30c",
   8856 => x"30c30c",
   8857 => x"30c30c",
   8858 => x"30c30c",
   8859 => x"30c30c",
   8860 => x"30c30c",
   8861 => x"30c30c",
   8862 => x"30c30c",
   8863 => x"30c30c",
   8864 => x"30c76e",
   8865 => x"ffffff",
   8866 => x"ffffff",
   8867 => x"ffffff",
   8868 => x"ffffff",
   8869 => x"ffffff",
   8870 => x"ffffff",
   8871 => x"ffffff",
   8872 => x"ffffff",
   8873 => x"ffffff",
   8874 => x"ffffff",
   8875 => x"ffffff",
   8876 => x"ffffff",
   8877 => x"ffffff",
   8878 => x"ffffff",
   8879 => x"ffffff",
   8880 => x"ffffff",
   8881 => x"ffffff",
   8882 => x"ffffff",
   8883 => x"ffffff",
   8884 => x"ffffff",
   8885 => x"ffffff",
   8886 => x"ffffff",
   8887 => x"ffffff",
   8888 => x"ffffff",
   8889 => x"ffffff",
   8890 => x"ffffff",
   8891 => x"ffffff",
   8892 => x"ffffff",
   8893 => x"ffffff",
   8894 => x"ffffff",
   8895 => x"ffffff",
   8896 => x"ffffff",
   8897 => x"ffffea",
   8898 => x"56afff",
   8899 => x"ffffff",
   8900 => x"ffffff",
   8901 => x"ffffff",
   8902 => x"ffffff",
   8903 => x"ffffff",
   8904 => x"ffffff",
   8905 => x"ffffff",
   8906 => x"ffffff",
   8907 => x"ffffff",
   8908 => x"ffffff",
   8909 => x"ffffff",
   8910 => x"ffffff",
   8911 => x"ffffff",
   8912 => x"ffffff",
   8913 => x"ffffff",
   8914 => x"ffffff",
   8915 => x"ffffff",
   8916 => x"ffffff",
   8917 => x"ffffff",
   8918 => x"ffffff",
   8919 => x"ffffff",
   8920 => x"ffffff",
   8921 => x"ffffff",
   8922 => x"ffffff",
   8923 => x"ffffff",
   8924 => x"ffffff",
   8925 => x"ffffff",
   8926 => x"ffffff",
   8927 => x"ffffff",
   8928 => x"ffffff",
   8929 => x"ffffff",
   8930 => x"ffffff",
   8931 => x"ffffff",
   8932 => x"ffffff",
   8933 => x"ffffff",
   8934 => x"ffffff",
   8935 => x"ffffff",
   8936 => x"ffffff",
   8937 => x"ffffff",
   8938 => x"ffffff",
   8939 => x"ffffff",
   8940 => x"ffffff",
   8941 => x"ffffff",
   8942 => x"ffffff",
   8943 => x"ffffff",
   8944 => x"ffffff",
   8945 => x"ffffff",
   8946 => x"ffffff",
   8947 => x"ffffff",
   8948 => x"ffffff",
   8949 => x"ffffff",
   8950 => x"ffffff",
   8951 => x"ffffff",
   8952 => x"ffffff",
   8953 => x"ffffff",
   8954 => x"ffffff",
   8955 => x"ffffff",
   8956 => x"ffffff",
   8957 => x"ffffff",
   8958 => x"ffffff",
   8959 => x"ffffff",
   8960 => x"ffffff",
   8961 => x"ffffff",
   8962 => x"ffffff",
   8963 => x"fffeb0",
   8964 => x"c30c30",
   8965 => x"c30c30",
   8966 => x"c30c30",
   8967 => x"c30c30",
   8968 => x"c30c30",
   8969 => x"c30c30",
   8970 => x"c30c30",
   8971 => x"c30c30",
   8972 => x"c30c30",
   8973 => x"c30c30",
   8974 => x"c30c30",
   8975 => x"c30c30",
   8976 => x"c30c30",
   8977 => x"c30c30",
   8978 => x"c30c30",
   8979 => x"c30c30",
   8980 => x"c30c30",
   8981 => x"c30c30",
   8982 => x"c30c30",
   8983 => x"c30c30",
   8984 => x"c30c30",
   8985 => x"c3063c",
   8986 => x"f3cf3c",
   8987 => x"f3cf3c",
   8988 => x"f3cf3c",
   8989 => x"f3cf3c",
   8990 => x"f3cf3c",
   8991 => x"f3cf3c",
   8992 => x"f3cf3c",
   8993 => x"f3cf3c",
   8994 => x"f3cf3c",
   8995 => x"f3cf3c",
   8996 => x"f3cf3c",
   8997 => x"f3cf3c",
   8998 => x"f3cf3c",
   8999 => x"f3cf3c",
   9000 => x"f3cf3c",
   9001 => x"f3cf3c",
   9002 => x"f3cf2c",
   9003 => x"30c30c",
   9004 => x"30c30c",
   9005 => x"30c30c",
   9006 => x"30c30c",
   9007 => x"30c30c",
   9008 => x"30c30c",
   9009 => x"30c30c",
   9010 => x"30c30c",
   9011 => x"30c30c",
   9012 => x"30c30c",
   9013 => x"30c30c",
   9014 => x"30c30c",
   9015 => x"30c30c",
   9016 => x"30c30c",
   9017 => x"30c30c",
   9018 => x"30c30c",
   9019 => x"30c30c",
   9020 => x"30c30c",
   9021 => x"30c30c",
   9022 => x"30c30c",
   9023 => x"30c30c",
   9024 => x"30c31d",
   9025 => x"ffffff",
   9026 => x"ffffff",
   9027 => x"ffffff",
   9028 => x"ffffff",
   9029 => x"ffffff",
   9030 => x"ffffff",
   9031 => x"ffffff",
   9032 => x"ffffff",
   9033 => x"ffffff",
   9034 => x"ffffff",
   9035 => x"ffffff",
   9036 => x"ffffff",
   9037 => x"ffffff",
   9038 => x"ffffff",
   9039 => x"ffffff",
   9040 => x"ffffff",
   9041 => x"ffffff",
   9042 => x"ffffff",
   9043 => x"ffffff",
   9044 => x"ffffff",
   9045 => x"ffffff",
   9046 => x"ffffff",
   9047 => x"ffffff",
   9048 => x"ffffff",
   9049 => x"ffffff",
   9050 => x"ffffff",
   9051 => x"ffffff",
   9052 => x"ffffff",
   9053 => x"ffffff",
   9054 => x"ffffff",
   9055 => x"ffffff",
   9056 => x"ffffff",
   9057 => x"fffa95",
   9058 => x"abffff",
   9059 => x"ffffff",
   9060 => x"ffffff",
   9061 => x"ffffff",
   9062 => x"ffffff",
   9063 => x"ffffff",
   9064 => x"ffffff",
   9065 => x"ffffff",
   9066 => x"ffffff",
   9067 => x"ffffff",
   9068 => x"ffffff",
   9069 => x"ffffff",
   9070 => x"ffffff",
   9071 => x"ffffff",
   9072 => x"ffffff",
   9073 => x"ffffff",
   9074 => x"ffffff",
   9075 => x"ffffff",
   9076 => x"ffffff",
   9077 => x"ffffff",
   9078 => x"ffffff",
   9079 => x"ffffff",
   9080 => x"ffffff",
   9081 => x"ffffff",
   9082 => x"ffffff",
   9083 => x"ffffff",
   9084 => x"ffffff",
   9085 => x"ffffff",
   9086 => x"ffffff",
   9087 => x"ffffff",
   9088 => x"ffffff",
   9089 => x"ffffff",
   9090 => x"ffffff",
   9091 => x"ffffff",
   9092 => x"ffffff",
   9093 => x"ffffff",
   9094 => x"ffffff",
   9095 => x"ffffff",
   9096 => x"ffffff",
   9097 => x"ffffff",
   9098 => x"ffffff",
   9099 => x"ffffff",
   9100 => x"ffffff",
   9101 => x"ffffff",
   9102 => x"ffffff",
   9103 => x"ffffff",
   9104 => x"ffffff",
   9105 => x"ffffff",
   9106 => x"ffffff",
   9107 => x"ffffff",
   9108 => x"ffffff",
   9109 => x"ffffff",
   9110 => x"ffffff",
   9111 => x"ffffff",
   9112 => x"ffffff",
   9113 => x"ffffff",
   9114 => x"ffffff",
   9115 => x"ffffff",
   9116 => x"ffffff",
   9117 => x"ffffff",
   9118 => x"ffffff",
   9119 => x"ffffff",
   9120 => x"ffffff",
   9121 => x"ffffff",
   9122 => x"ffffff",
   9123 => x"fffd70",
   9124 => x"c30c30",
   9125 => x"c30c30",
   9126 => x"c30c30",
   9127 => x"c30c30",
   9128 => x"c30c30",
   9129 => x"c30c30",
   9130 => x"c30c30",
   9131 => x"c30c30",
   9132 => x"c30c30",
   9133 => x"c30c30",
   9134 => x"c30c30",
   9135 => x"c30c30",
   9136 => x"c30c30",
   9137 => x"c30c30",
   9138 => x"c30c30",
   9139 => x"c30c30",
   9140 => x"c30c30",
   9141 => x"c30c30",
   9142 => x"c30c30",
   9143 => x"c30c30",
   9144 => x"c30c30",
   9145 => x"c24b3c",
   9146 => x"f3cf3c",
   9147 => x"f3cf3c",
   9148 => x"f3cf3c",
   9149 => x"f3cf3c",
   9150 => x"f3cf3c",
   9151 => x"f3cf3c",
   9152 => x"f3cf3c",
   9153 => x"f3cf3c",
   9154 => x"f3cf3c",
   9155 => x"f3cf3c",
   9156 => x"f3cf3c",
   9157 => x"f3cf3c",
   9158 => x"f3cf3c",
   9159 => x"f3cf3c",
   9160 => x"f3cf3c",
   9161 => x"f3cf3c",
   9162 => x"f3cf3c",
   9163 => x"70c30c",
   9164 => x"30c30c",
   9165 => x"30c30c",
   9166 => x"30c30c",
   9167 => x"30c30c",
   9168 => x"30c30c",
   9169 => x"30c30c",
   9170 => x"30c30c",
   9171 => x"30c30c",
   9172 => x"30c30c",
   9173 => x"30c30c",
   9174 => x"30c30c",
   9175 => x"30c30c",
   9176 => x"30c30c",
   9177 => x"30c30c",
   9178 => x"30c30c",
   9179 => x"30c30c",
   9180 => x"30c30c",
   9181 => x"30c30c",
   9182 => x"30c30c",
   9183 => x"30c30c",
   9184 => x"30c30c",
   9185 => x"bbffff",
   9186 => x"ffffff",
   9187 => x"ffffff",
   9188 => x"ffffff",
   9189 => x"ffffff",
   9190 => x"ffffff",
   9191 => x"ffffff",
   9192 => x"ffffff",
   9193 => x"ffffff",
   9194 => x"ffffff",
   9195 => x"ffffff",
   9196 => x"ffffff",
   9197 => x"ffffff",
   9198 => x"ffffff",
   9199 => x"ffffff",
   9200 => x"ffffff",
   9201 => x"ffffff",
   9202 => x"ffffff",
   9203 => x"ffffff",
   9204 => x"ffffff",
   9205 => x"ffffff",
   9206 => x"ffffff",
   9207 => x"ffffff",
   9208 => x"ffffff",
   9209 => x"ffffff",
   9210 => x"ffffff",
   9211 => x"ffffff",
   9212 => x"ffffff",
   9213 => x"ffffff",
   9214 => x"ffffff",
   9215 => x"ffffff",
   9216 => x"ffffff",
   9217 => x"fea56a",
   9218 => x"ffffff",
   9219 => x"ffffff",
   9220 => x"ffffff",
   9221 => x"ffffff",
   9222 => x"ffffff",
   9223 => x"ffffff",
   9224 => x"ffffff",
   9225 => x"ffffff",
   9226 => x"ffffff",
   9227 => x"ffffff",
   9228 => x"ffffff",
   9229 => x"ffffff",
   9230 => x"ffffff",
   9231 => x"ffffff",
   9232 => x"ffffff",
   9233 => x"ffffff",
   9234 => x"ffffff",
   9235 => x"ffffff",
   9236 => x"ffffff",
   9237 => x"ffffff",
   9238 => x"ffffff",
   9239 => x"ffffff",
   9240 => x"ffffff",
   9241 => x"ffffff",
   9242 => x"ffffff",
   9243 => x"ffffff",
   9244 => x"ffffff",
   9245 => x"ffffff",
   9246 => x"ffffff",
   9247 => x"ffffff",
   9248 => x"ffffff",
   9249 => x"ffffff",
   9250 => x"ffffff",
   9251 => x"ffffff",
   9252 => x"ffffff",
   9253 => x"ffffff",
   9254 => x"ffffff",
   9255 => x"ffffff",
   9256 => x"ffffff",
   9257 => x"ffffff",
   9258 => x"ffffff",
   9259 => x"ffffff",
   9260 => x"ffffff",
   9261 => x"ffffff",
   9262 => x"ffffff",
   9263 => x"ffffff",
   9264 => x"ffffff",
   9265 => x"ffffff",
   9266 => x"ffffff",
   9267 => x"ffffff",
   9268 => x"ffffff",
   9269 => x"ffffff",
   9270 => x"ffffff",
   9271 => x"ffffff",
   9272 => x"ffffff",
   9273 => x"ffffff",
   9274 => x"ffffff",
   9275 => x"ffffff",
   9276 => x"ffffff",
   9277 => x"ffffff",
   9278 => x"ffffff",
   9279 => x"ffffff",
   9280 => x"ffffff",
   9281 => x"ffffff",
   9282 => x"ffffff",
   9283 => x"ffac30",
   9284 => x"c30c30",
   9285 => x"c30c30",
   9286 => x"c30c30",
   9287 => x"c30c30",
   9288 => x"c30c30",
   9289 => x"c30c30",
   9290 => x"c30c30",
   9291 => x"c30c30",
   9292 => x"c30c30",
   9293 => x"c30c30",
   9294 => x"c30c30",
   9295 => x"c30c30",
   9296 => x"c30c30",
   9297 => x"c30c30",
   9298 => x"c30c30",
   9299 => x"c30c30",
   9300 => x"c30c30",
   9301 => x"c30c30",
   9302 => x"c30c30",
   9303 => x"c30c30",
   9304 => x"c30c30",
   9305 => x"92cf3c",
   9306 => x"f3cf3c",
   9307 => x"f3cf3c",
   9308 => x"f3cf3c",
   9309 => x"f3cf3c",
   9310 => x"f3cf3c",
   9311 => x"f3cf3c",
   9312 => x"f3cf3c",
   9313 => x"f3cf3c",
   9314 => x"f3cf3c",
   9315 => x"f3cf3c",
   9316 => x"f3cf3c",
   9317 => x"f3cf3c",
   9318 => x"f3cf3c",
   9319 => x"f3cf3c",
   9320 => x"f3cf3c",
   9321 => x"f3cf3c",
   9322 => x"f3cf3c",
   9323 => x"b1c30c",
   9324 => x"30c30c",
   9325 => x"30c30c",
   9326 => x"30c30c",
   9327 => x"30c30c",
   9328 => x"30c30c",
   9329 => x"30c30c",
   9330 => x"30c30c",
   9331 => x"30c30c",
   9332 => x"30c30c",
   9333 => x"30c30c",
   9334 => x"30c30c",
   9335 => x"30c30c",
   9336 => x"30c30c",
   9337 => x"30c30c",
   9338 => x"30c30c",
   9339 => x"30c30c",
   9340 => x"30c30c",
   9341 => x"30c30c",
   9342 => x"30c30c",
   9343 => x"30c30c",
   9344 => x"30c30c",
   9345 => x"76efff",
   9346 => x"ffffff",
   9347 => x"ffffff",
   9348 => x"ffffff",
   9349 => x"ffffff",
   9350 => x"ffffff",
   9351 => x"ffffff",
   9352 => x"ffffff",
   9353 => x"ffffff",
   9354 => x"ffffff",
   9355 => x"ffffff",
   9356 => x"ffffff",
   9357 => x"ffffff",
   9358 => x"ffffff",
   9359 => x"ffffff",
   9360 => x"ffffff",
   9361 => x"ffffff",
   9362 => x"ffffff",
   9363 => x"ffffff",
   9364 => x"ffffff",
   9365 => x"ffffff",
   9366 => x"ffffff",
   9367 => x"ffffff",
   9368 => x"ffffff",
   9369 => x"ffffff",
   9370 => x"ffffff",
   9371 => x"ffffff",
   9372 => x"ffffff",
   9373 => x"ffffff",
   9374 => x"ffffff",
   9375 => x"ffffff",
   9376 => x"ffffff",
   9377 => x"a95abf",
   9378 => x"ffffff",
   9379 => x"ffffff",
   9380 => x"ffffff",
   9381 => x"ffffff",
   9382 => x"ffffff",
   9383 => x"ffffff",
   9384 => x"ffffff",
   9385 => x"ffffff",
   9386 => x"ffffff",
   9387 => x"ffffff",
   9388 => x"ffffff",
   9389 => x"ffffff",
   9390 => x"ffffff",
   9391 => x"ffffff",
   9392 => x"ffffff",
   9393 => x"ffffff",
   9394 => x"ffffff",
   9395 => x"ffffff",
   9396 => x"ffffff",
   9397 => x"ffffff",
   9398 => x"ffffff",
   9399 => x"ffffff",
   9400 => x"ffffff",
   9401 => x"ffffff",
   9402 => x"ffffff",
   9403 => x"ffffff",
   9404 => x"ffffff",
   9405 => x"ffffff",
   9406 => x"ffffff",
   9407 => x"ffffff",
   9408 => x"ffffff",
   9409 => x"ffffff",
   9410 => x"ffffff",
   9411 => x"ffffff",
   9412 => x"ffffff",
   9413 => x"ffffff",
   9414 => x"ffffff",
   9415 => x"ffffff",
   9416 => x"ffffff",
   9417 => x"ffffff",
   9418 => x"ffffff",
   9419 => x"ffffff",
   9420 => x"ffffff",
   9421 => x"ffffff",
   9422 => x"ffffff",
   9423 => x"ffffff",
   9424 => x"ffffff",
   9425 => x"ffffff",
   9426 => x"ffffff",
   9427 => x"ffffff",
   9428 => x"ffffff",
   9429 => x"ffffff",
   9430 => x"ffffff",
   9431 => x"ffffff",
   9432 => x"ffffff",
   9433 => x"ffffff",
   9434 => x"ffffff",
   9435 => x"ffffff",
   9436 => x"ffffff",
   9437 => x"ffffff",
   9438 => x"ffffff",
   9439 => x"ffffff",
   9440 => x"ffffff",
   9441 => x"ffffff",
   9442 => x"ffffff",
   9443 => x"eb5c30",
   9444 => x"c30c30",
   9445 => x"c30c30",
   9446 => x"c30c30",
   9447 => x"c30c30",
   9448 => x"c30c30",
   9449 => x"c30c30",
   9450 => x"c30c30",
   9451 => x"c30c30",
   9452 => x"c30c30",
   9453 => x"c30c30",
   9454 => x"c30c30",
   9455 => x"c30c30",
   9456 => x"c30c30",
   9457 => x"c30c30",
   9458 => x"c30c30",
   9459 => x"c30c30",
   9460 => x"c30c30",
   9461 => x"c30c30",
   9462 => x"c30c30",
   9463 => x"c30c30",
   9464 => x"c30c30",
   9465 => x"a3cf3c",
   9466 => x"f3cf3c",
   9467 => x"f3cf3c",
   9468 => x"f3cf3c",
   9469 => x"f3cf3c",
   9470 => x"f3cf3c",
   9471 => x"f3cf3c",
   9472 => x"f3cf3c",
   9473 => x"f3cf3c",
   9474 => x"f3cf3c",
   9475 => x"f3cf3c",
   9476 => x"f3cf3c",
   9477 => x"f3cf3c",
   9478 => x"f3cf3c",
   9479 => x"f3cf3c",
   9480 => x"f3cf3c",
   9481 => x"f3cf3c",
   9482 => x"f3cf3c",
   9483 => x"f2c30c",
   9484 => x"30c30c",
   9485 => x"30c30c",
   9486 => x"30c30c",
   9487 => x"30c30c",
   9488 => x"30c30c",
   9489 => x"30c30c",
   9490 => x"30c30c",
   9491 => x"30c30c",
   9492 => x"30c30c",
   9493 => x"30c30c",
   9494 => x"30c30c",
   9495 => x"30c30c",
   9496 => x"30c30c",
   9497 => x"30c30c",
   9498 => x"30c30c",
   9499 => x"30c30c",
   9500 => x"30c30c",
   9501 => x"30c30c",
   9502 => x"30c30c",
   9503 => x"30c30c",
   9504 => x"30c30c",
   9505 => x"31dfff",
   9506 => x"ffffff",
   9507 => x"ffffff",
   9508 => x"ffffff",
   9509 => x"ffffff",
   9510 => x"ffffff",
   9511 => x"ffffff",
   9512 => x"ffffff",
   9513 => x"ffffff",
   9514 => x"ffffff",
   9515 => x"ffffff",
   9516 => x"ffffff",
   9517 => x"ffffff",
   9518 => x"ffffff",
   9519 => x"ffffff",
   9520 => x"ffffff",
   9521 => x"ffffff",
   9522 => x"ffffff",
   9523 => x"ffffff",
   9524 => x"ffffff",
   9525 => x"ffffff",
   9526 => x"ffffff",
   9527 => x"ffffff",
   9528 => x"ffffff",
   9529 => x"ffffff",
   9530 => x"ffffff",
   9531 => x"ffffff",
   9532 => x"ffffff",
   9533 => x"ffffff",
   9534 => x"ffffff",
   9535 => x"ffffff",
   9536 => x"ffffea",
   9537 => x"56afff",
   9538 => x"ffffff",
   9539 => x"ffffff",
   9540 => x"ffffff",
   9541 => x"ffffff",
   9542 => x"ffffff",
   9543 => x"ffffff",
   9544 => x"ffffff",
   9545 => x"ffffff",
   9546 => x"ffffff",
   9547 => x"ffffff",
   9548 => x"ffffff",
   9549 => x"ffffff",
   9550 => x"ffffff",
   9551 => x"ffffff",
   9552 => x"ffffff",
   9553 => x"ffffff",
   9554 => x"ffffff",
   9555 => x"ffffff",
   9556 => x"ffffff",
   9557 => x"ffffff",
   9558 => x"ffffff",
   9559 => x"ffffff",
   9560 => x"ffffff",
   9561 => x"ffffff",
   9562 => x"ffffff",
   9563 => x"ffffff",
   9564 => x"ffffff",
   9565 => x"ffffff",
   9566 => x"ffffff",
   9567 => x"ffffff",
   9568 => x"ffffff",
   9569 => x"ffffff",
   9570 => x"ffffff",
   9571 => x"ffffff",
   9572 => x"ffffff",
   9573 => x"ffffff",
   9574 => x"ffffff",
   9575 => x"ffffff",
   9576 => x"ffffff",
   9577 => x"ffffff",
   9578 => x"ffffff",
   9579 => x"ffffff",
   9580 => x"ffffff",
   9581 => x"ffffff",
   9582 => x"ffffff",
   9583 => x"ffffff",
   9584 => x"ffffff",
   9585 => x"ffffff",
   9586 => x"ffffff",
   9587 => x"ffffff",
   9588 => x"ffffff",
   9589 => x"ffffff",
   9590 => x"ffffff",
   9591 => x"ffffff",
   9592 => x"ffffff",
   9593 => x"ffffff",
   9594 => x"ffffff",
   9595 => x"ffffff",
   9596 => x"ffffff",
   9597 => x"ffffff",
   9598 => x"ffffff",
   9599 => x"ffffff",
   9600 => x"ffffff",
   9601 => x"ffffff",
   9602 => x"ffffff",
   9603 => x"d70c30",
   9604 => x"c30c30",
   9605 => x"c30c30",
   9606 => x"c30c30",
   9607 => x"c30c30",
   9608 => x"c30c30",
   9609 => x"c30c30",
   9610 => x"c30c30",
   9611 => x"c30c30",
   9612 => x"c30c30",
   9613 => x"c30c30",
   9614 => x"c30c30",
   9615 => x"c30c30",
   9616 => x"c30c30",
   9617 => x"c30c30",
   9618 => x"c30c30",
   9619 => x"c30c30",
   9620 => x"c30c30",
   9621 => x"c30c30",
   9622 => x"c30c30",
   9623 => x"c30c30",
   9624 => x"c30c24",
   9625 => x"b3cf3c",
   9626 => x"f3cf3c",
   9627 => x"f3cf3c",
   9628 => x"f3cf3c",
   9629 => x"f3cf3c",
   9630 => x"f3cf3c",
   9631 => x"f3cf3c",
   9632 => x"f3cf3c",
   9633 => x"f3cf3c",
   9634 => x"f3cf3c",
   9635 => x"f3cf3c",
   9636 => x"f3cf3c",
   9637 => x"f3cf3c",
   9638 => x"f3cf3c",
   9639 => x"f3cf3c",
   9640 => x"f3cf3c",
   9641 => x"f3cf3c",
   9642 => x"f3cf3c",
   9643 => x"f3c70c",
   9644 => x"30c30c",
   9645 => x"30c30c",
   9646 => x"30c30c",
   9647 => x"30c30c",
   9648 => x"30c30c",
   9649 => x"30c30c",
   9650 => x"30c30c",
   9651 => x"30c30c",
   9652 => x"30c30c",
   9653 => x"30c30c",
   9654 => x"30c30c",
   9655 => x"30c30c",
   9656 => x"30c30c",
   9657 => x"30c30c",
   9658 => x"30c30c",
   9659 => x"30c30c",
   9660 => x"30c30c",
   9661 => x"30c30c",
   9662 => x"30c30c",
   9663 => x"30c30c",
   9664 => x"30c30c",
   9665 => x"30cbbf",
   9666 => x"ffffff",
   9667 => x"ffffff",
   9668 => x"ffffff",
   9669 => x"ffffff",
   9670 => x"ffffff",
   9671 => x"ffffff",
   9672 => x"ffffff",
   9673 => x"ffffff",
   9674 => x"ffffff",
   9675 => x"ffffff",
   9676 => x"ffffff",
   9677 => x"ffffff",
   9678 => x"ffffff",
   9679 => x"ffffff",
   9680 => x"ffffff",
   9681 => x"ffffff",
   9682 => x"ffffff",
   9683 => x"ffffff",
   9684 => x"ffffff",
   9685 => x"ffffff",
   9686 => x"ffffff",
   9687 => x"ffffff",
   9688 => x"ffffff",
   9689 => x"ffffff",
   9690 => x"ffffff",
   9691 => x"ffffff",
   9692 => x"ffffff",
   9693 => x"ffffff",
   9694 => x"ffffff",
   9695 => x"ffffff",
   9696 => x"fffa95",
   9697 => x"abffff",
   9698 => x"ffffff",
   9699 => x"ffffff",
   9700 => x"ffffff",
   9701 => x"ffffff",
   9702 => x"ffffff",
   9703 => x"ffffff",
   9704 => x"ffffff",
   9705 => x"ffffff",
   9706 => x"ffffff",
   9707 => x"ffffff",
   9708 => x"ffffff",
   9709 => x"ffffff",
   9710 => x"ffffff",
   9711 => x"ffffff",
   9712 => x"ffffff",
   9713 => x"ffffff",
   9714 => x"ffffff",
   9715 => x"ffffff",
   9716 => x"ffffff",
   9717 => x"ffffff",
   9718 => x"ffffff",
   9719 => x"ffffff",
   9720 => x"ffffff",
   9721 => x"ffffff",
   9722 => x"ffffff",
   9723 => x"ffffff",
   9724 => x"ffffff",
   9725 => x"ffffff",
   9726 => x"ffffff",
   9727 => x"ffffff",
   9728 => x"ffffff",
   9729 => x"ffffff",
   9730 => x"ffffff",
   9731 => x"ffffff",
   9732 => x"ffffff",
   9733 => x"ffffff",
   9734 => x"ffffff",
   9735 => x"ffffff",
   9736 => x"ffffff",
   9737 => x"ffffff",
   9738 => x"ffffff",
   9739 => x"ffffff",
   9740 => x"ffffff",
   9741 => x"ffffff",
   9742 => x"ffffff",
   9743 => x"ffffff",
   9744 => x"ffffff",
   9745 => x"ffffff",
   9746 => x"ffffff",
   9747 => x"ffffff",
   9748 => x"ffffff",
   9749 => x"ffffff",
   9750 => x"ffffff",
   9751 => x"ffffff",
   9752 => x"ffffff",
   9753 => x"ffffff",
   9754 => x"ffffff",
   9755 => x"ffffff",
   9756 => x"ffffff",
   9757 => x"ffffff",
   9758 => x"ffffff",
   9759 => x"ffffff",
   9760 => x"ffffff",
   9761 => x"ffffff",
   9762 => x"fffffa",
   9763 => x"d70c30",
   9764 => x"c30c30",
   9765 => x"c30c30",
   9766 => x"c30c30",
   9767 => x"c30c30",
   9768 => x"c30c30",
   9769 => x"c30c30",
   9770 => x"c30c30",
   9771 => x"c30c30",
   9772 => x"c30c30",
   9773 => x"c30c30",
   9774 => x"c30c30",
   9775 => x"c30c30",
   9776 => x"c30c30",
   9777 => x"c30c30",
   9778 => x"c30c30",
   9779 => x"c30c30",
   9780 => x"c30c30",
   9781 => x"c30c30",
   9782 => x"c30c30",
   9783 => x"c30c30",
   9784 => x"c30c28",
   9785 => x"f3cf3c",
   9786 => x"f3cf3c",
   9787 => x"f3cf3c",
   9788 => x"f3cf3c",
   9789 => x"f3cf3c",
   9790 => x"f3cf3c",
   9791 => x"f3cf3c",
   9792 => x"f3cf3c",
   9793 => x"f3cf3c",
   9794 => x"f3cf3c",
   9795 => x"f3cf3c",
   9796 => x"f3cf3c",
   9797 => x"f3cf3c",
   9798 => x"f3cf3c",
   9799 => x"f3cf3c",
   9800 => x"f3cf3c",
   9801 => x"f3cf3c",
   9802 => x"f3cf3c",
   9803 => x"f3cb0c",
   9804 => x"30c30c",
   9805 => x"30c30c",
   9806 => x"30c30c",
   9807 => x"30c30c",
   9808 => x"30c30c",
   9809 => x"30c30c",
   9810 => x"30c30c",
   9811 => x"30c30c",
   9812 => x"30c30c",
   9813 => x"30c30c",
   9814 => x"30c30c",
   9815 => x"30c30c",
   9816 => x"30c30c",
   9817 => x"30c30c",
   9818 => x"30c30c",
   9819 => x"30c30c",
   9820 => x"30c30c",
   9821 => x"30c30c",
   9822 => x"30c30c",
   9823 => x"30c30c",
   9824 => x"30c30c",
   9825 => x"30c77f",
   9826 => x"ffffff",
   9827 => x"ffffff",
   9828 => x"ffffff",
   9829 => x"ffffff",
   9830 => x"ffffff",
   9831 => x"ffffff",
   9832 => x"ffffff",
   9833 => x"ffffff",
   9834 => x"ffffff",
   9835 => x"ffffff",
   9836 => x"ffffff",
   9837 => x"ffffff",
   9838 => x"ffffff",
   9839 => x"ffffff",
   9840 => x"ffffff",
   9841 => x"ffffff",
   9842 => x"ffffff",
   9843 => x"ffffff",
   9844 => x"ffffff",
   9845 => x"ffffff",
   9846 => x"ffffff",
   9847 => x"ffffff",
   9848 => x"ffffff",
   9849 => x"ffffff",
   9850 => x"ffffff",
   9851 => x"ffffff",
   9852 => x"ffffff",
   9853 => x"ffffff",
   9854 => x"ffffff",
   9855 => x"ffffff",
   9856 => x"fea56a",
   9857 => x"ffffff",
   9858 => x"ffffff",
   9859 => x"ffffff",
   9860 => x"ffffff",
   9861 => x"ffffff",
   9862 => x"ffffff",
   9863 => x"ffffff",
   9864 => x"ffffff",
   9865 => x"ffffff",
   9866 => x"ffffff",
   9867 => x"ffffff",
   9868 => x"ffffff",
   9869 => x"ffffff",
   9870 => x"ffffff",
   9871 => x"ffffff",
   9872 => x"ffffff",
   9873 => x"ffffff",
   9874 => x"ffffff",
   9875 => x"ffffff",
   9876 => x"ffffff",
   9877 => x"ffffff",
   9878 => x"ffffff",
   9879 => x"ffffff",
   9880 => x"ffffff",
   9881 => x"ffffff",
   9882 => x"ffffff",
   9883 => x"ffffff",
   9884 => x"ffffff",
   9885 => x"ffffff",
   9886 => x"ffffff",
   9887 => x"ffffff",
   9888 => x"ffffff",
   9889 => x"ffffff",
   9890 => x"ffffff",
   9891 => x"ffffff",
   9892 => x"ffffff",
   9893 => x"ffffff",
   9894 => x"ffffff",
   9895 => x"ffffff",
   9896 => x"ffffff",
   9897 => x"ffffff",
   9898 => x"ffffff",
   9899 => x"ffffff",
   9900 => x"ffffff",
   9901 => x"ffffff",
   9902 => x"ffffff",
   9903 => x"ffffff",
   9904 => x"ffffff",
   9905 => x"ffffff",
   9906 => x"ffffff",
   9907 => x"ffffff",
   9908 => x"ffffff",
   9909 => x"ffffff",
   9910 => x"ffffff",
   9911 => x"ffffff",
   9912 => x"ffffff",
   9913 => x"ffffff",
   9914 => x"ffffff",
   9915 => x"ffffff",
   9916 => x"ffffff",
   9917 => x"ffffff",
   9918 => x"ffffff",
   9919 => x"ffffff",
   9920 => x"ffffff",
   9921 => x"ffffff",
   9922 => x"fffff5",
   9923 => x"c30c30",
   9924 => x"c30c30",
   9925 => x"c30c30",
   9926 => x"c30c30",
   9927 => x"c30c30",
   9928 => x"c30c30",
   9929 => x"c30c30",
   9930 => x"c30c30",
   9931 => x"c30c30",
   9932 => x"c30c30",
   9933 => x"c30c30",
   9934 => x"c30c30",
   9935 => x"c30c30",
   9936 => x"c30c30",
   9937 => x"c30c30",
   9938 => x"c30c30",
   9939 => x"c30c30",
   9940 => x"c30c30",
   9941 => x"c30c30",
   9942 => x"c30c30",
   9943 => x"c30c30",
   9944 => x"c3092c",
   9945 => x"f3cf3c",
   9946 => x"f3cf3c",
   9947 => x"f3cf3c",
   9948 => x"f3cf3c",
   9949 => x"f3cf3c",
   9950 => x"f3cf3c",
   9951 => x"f3cf3c",
   9952 => x"f3cf3c",
   9953 => x"f3cf3c",
   9954 => x"f3cf3c",
   9955 => x"f3cf3c",
   9956 => x"f3cf3c",
   9957 => x"f3cf3c",
   9958 => x"f3cf3c",
   9959 => x"f3cf3c",
   9960 => x"f3cf3c",
   9961 => x"f3cf3c",
   9962 => x"f3cf3c",
   9963 => x"f3cf1c",
   9964 => x"30c30c",
   9965 => x"30c30c",
   9966 => x"30c30c",
   9967 => x"30c30c",
   9968 => x"30c30c",
   9969 => x"30c30c",
   9970 => x"30c30c",
   9971 => x"30c30c",
   9972 => x"30c30c",
   9973 => x"30c30c",
   9974 => x"30c30c",
   9975 => x"30c30c",
   9976 => x"30c30c",
   9977 => x"30c30c",
   9978 => x"30c30c",
   9979 => x"30c30c",
   9980 => x"30c30c",
   9981 => x"30c30c",
   9982 => x"30c30c",
   9983 => x"30c30c",
   9984 => x"30c30c",
   9985 => x"30c32e",
   9986 => x"ffffff",
   9987 => x"ffffff",
   9988 => x"ffffff",
   9989 => x"ffffff",
   9990 => x"ffffff",
   9991 => x"ffffff",
   9992 => x"ffffff",
   9993 => x"ffffff",
   9994 => x"ffffff",
   9995 => x"ffffff",
   9996 => x"ffffff",
   9997 => x"ffffff",
   9998 => x"ffffff",
   9999 => x"ffffff",
   10000 => x"ffffff",
   10001 => x"ffffff",
   10002 => x"ffffff",
   10003 => x"ffffff",
   10004 => x"ffffff",
   10005 => x"ffffff",
   10006 => x"ffffff",
   10007 => x"ffffff",
   10008 => x"ffffff",
   10009 => x"ffffff",
   10010 => x"ffffff",
   10011 => x"ffffff",
   10012 => x"ffffff",
   10013 => x"ffffff",
   10014 => x"ffffff",
   10015 => x"ffffff",
   10016 => x"a95abf",
   10017 => x"ffffff",
   10018 => x"ffffff",
   10019 => x"ffffff",
   10020 => x"ffffff",
   10021 => x"ffffff",
   10022 => x"ffffff",
   10023 => x"ffffff",
   10024 => x"ffffff",
   10025 => x"ffffff",
   10026 => x"ffffff",
   10027 => x"ffffff",
   10028 => x"ffffff",
   10029 => x"ffffff",
   10030 => x"ffffff",
   10031 => x"ffffff",
   10032 => x"ffffff",
   10033 => x"ffffff",
   10034 => x"ffffff",
   10035 => x"ffffff",
   10036 => x"ffffff",
   10037 => x"ffffff",
   10038 => x"ffffff",
   10039 => x"ffffff",
   10040 => x"ffffff",
   10041 => x"ffffff",
   10042 => x"ffffff",
   10043 => x"ffffff",
   10044 => x"ffffff",
   10045 => x"ffffff",
   10046 => x"ffffff",
   10047 => x"ffffff",
   10048 => x"ffffff",
   10049 => x"ffffff",
   10050 => x"ffffff",
   10051 => x"ffffff",
   10052 => x"ffffff",
   10053 => x"ffffff",
   10054 => x"ffffff",
   10055 => x"ffffff",
   10056 => x"ffffff",
   10057 => x"ffffff",
   10058 => x"ffffff",
   10059 => x"ffffff",
   10060 => x"ffffff",
   10061 => x"ffffff",
   10062 => x"ffffff",
   10063 => x"ffffff",
   10064 => x"ffffff",
   10065 => x"ffffff",
   10066 => x"ffffff",
   10067 => x"ffffff",
   10068 => x"ffffff",
   10069 => x"ffffff",
   10070 => x"ffffff",
   10071 => x"ffffff",
   10072 => x"ffffff",
   10073 => x"ffffff",
   10074 => x"ffffff",
   10075 => x"ffffff",
   10076 => x"ffffff",
   10077 => x"ffffff",
   10078 => x"ffffff",
   10079 => x"ffffff",
   10080 => x"ffffff",
   10081 => x"ffffff",
   10082 => x"fffeb5",
   10083 => x"c30c30",
   10084 => x"c30c30",
   10085 => x"c30c30",
   10086 => x"c30c30",
   10087 => x"c30c30",
   10088 => x"c30c30",
   10089 => x"c30c30",
   10090 => x"c30c30",
   10091 => x"c30c30",
   10092 => x"c30c30",
   10093 => x"c30c30",
   10094 => x"c30c30",
   10095 => x"c30c30",
   10096 => x"c30c30",
   10097 => x"c30c30",
   10098 => x"c30c30",
   10099 => x"c30c30",
   10100 => x"c30c30",
   10101 => x"c30c30",
   10102 => x"c30c30",
   10103 => x"c30c30",
   10104 => x"c30a3c",
   10105 => x"f3cf3c",
   10106 => x"f3cf3c",
   10107 => x"f3cf3c",
   10108 => x"f3cf3c",
   10109 => x"f3cf3c",
   10110 => x"f3cf3c",
   10111 => x"f3cf3c",
   10112 => x"f3cf3c",
   10113 => x"f3cf3c",
   10114 => x"f3cf3c",
   10115 => x"f3cf3c",
   10116 => x"f3cf3c",
   10117 => x"f3cf3c",
   10118 => x"f3cf3c",
   10119 => x"f3cf3c",
   10120 => x"f3cf3c",
   10121 => x"f3cf3c",
   10122 => x"f3cf3c",
   10123 => x"f3cf2c",
   10124 => x"30c30c",
   10125 => x"30c30c",
   10126 => x"30c30c",
   10127 => x"30c30c",
   10128 => x"30c30c",
   10129 => x"30c30c",
   10130 => x"30c30c",
   10131 => x"30c30c",
   10132 => x"30c30c",
   10133 => x"30c30c",
   10134 => x"30c30c",
   10135 => x"30c30c",
   10136 => x"30c30c",
   10137 => x"30c30c",
   10138 => x"30c30c",
   10139 => x"30c30c",
   10140 => x"30c30c",
   10141 => x"30c30c",
   10142 => x"30c30c",
   10143 => x"30c30c",
   10144 => x"30c30c",
   10145 => x"30c31d",
   10146 => x"ffffff",
   10147 => x"ffffff",
   10148 => x"ffffff",
   10149 => x"ffffff",
   10150 => x"ffffff",
   10151 => x"ffffff",
   10152 => x"ffffff",
   10153 => x"ffffff",
   10154 => x"ffffff",
   10155 => x"ffffff",
   10156 => x"ffffff",
   10157 => x"ffffff",
   10158 => x"ffffff",
   10159 => x"ffffff",
   10160 => x"ffffff",
   10161 => x"ffffff",
   10162 => x"ffffff",
   10163 => x"ffffff",
   10164 => x"ffffff",
   10165 => x"ffffff",
   10166 => x"ffffff",
   10167 => x"ffffff",
   10168 => x"ffffff",
   10169 => x"ffffff",
   10170 => x"ffffff",
   10171 => x"ffffff",
   10172 => x"ffffff",
   10173 => x"ffffff",
   10174 => x"ffffff",
   10175 => x"ffffea",
   10176 => x"56afff",
   10177 => x"ffffff",
   10178 => x"ffffff",
   10179 => x"ffffff",
   10180 => x"ffffff",
   10181 => x"ffffff",
   10182 => x"ffffff",
   10183 => x"ffffff",
   10184 => x"ffffff",
   10185 => x"ffffff",
   10186 => x"ffffff",
   10187 => x"ffffff",
   10188 => x"ffffff",
   10189 => x"ffffff",
   10190 => x"ffffff",
   10191 => x"ffffff",
   10192 => x"ffffff",
   10193 => x"ffffff",
   10194 => x"ffffff",
   10195 => x"ffffff",
   10196 => x"ffffff",
   10197 => x"ffffff",
   10198 => x"ffffff",
   10199 => x"ffffff",
   10200 => x"ffffff",
   10201 => x"ffffff",
   10202 => x"ffffff",
   10203 => x"ffffff",
   10204 => x"ffffff",
   10205 => x"ffffff",
   10206 => x"ffffff",
   10207 => x"ffffff",
   10208 => x"ffffff",
   10209 => x"ffffff",
   10210 => x"ffffff",
   10211 => x"ffffff",
   10212 => x"ffffff",
   10213 => x"ffffff",
   10214 => x"ffffff",
   10215 => x"ffffff",
   10216 => x"ffffff",
   10217 => x"ffffff",
   10218 => x"ffffff",
   10219 => x"ffffff",
   10220 => x"ffffff",
   10221 => x"ffffff",
   10222 => x"ffffff",
   10223 => x"ffffff",
   10224 => x"ffffff",
   10225 => x"ffffff",
   10226 => x"ffffff",
   10227 => x"ffffff",
   10228 => x"ffffff",
   10229 => x"ffffff",
   10230 => x"ffffff",
   10231 => x"ffffff",
   10232 => x"ffffff",
   10233 => x"ffffff",
   10234 => x"ffffff",
   10235 => x"ffffff",
   10236 => x"ffffff",
   10237 => x"ffffff",
   10238 => x"ffffff",
   10239 => x"ffffff",
   10240 => x"ffffff",
   10241 => x"ffffff",
   10242 => x"fffd70",
   10243 => x"c30c30",
   10244 => x"c30c30",
   10245 => x"c30c30",
   10246 => x"c30c30",
   10247 => x"c30c30",
   10248 => x"c30c30",
   10249 => x"c30c30",
   10250 => x"c30c30",
   10251 => x"c30c30",
   10252 => x"c30c30",
   10253 => x"c30c30",
   10254 => x"c30c30",
   10255 => x"c30c30",
   10256 => x"c30c30",
   10257 => x"c30c30",
   10258 => x"c30c30",
   10259 => x"c30c30",
   10260 => x"c30c30",
   10261 => x"c30c30",
   10262 => x"c30c30",
   10263 => x"c30c30",
   10264 => x"c24b3c",
   10265 => x"f3cf3c",
   10266 => x"f3cf3c",
   10267 => x"f3cf3c",
   10268 => x"f3cf3c",
   10269 => x"f3cf3c",
   10270 => x"f3cf3c",
   10271 => x"f3cf3c",
   10272 => x"f3cf3c",
   10273 => x"f3cf3c",
   10274 => x"f3cf3c",
   10275 => x"f3cf3c",
   10276 => x"f3cf3c",
   10277 => x"f3cf3c",
   10278 => x"f3cf3c",
   10279 => x"f3cf3c",
   10280 => x"f3cf3c",
   10281 => x"f3cf3c",
   10282 => x"f3cf3c",
   10283 => x"f3cf2c",
   10284 => x"70c30c",
   10285 => x"30c30c",
   10286 => x"30c30c",
   10287 => x"30c30c",
   10288 => x"30c30c",
   10289 => x"30c30c",
   10290 => x"30c30c",
   10291 => x"30c30c",
   10292 => x"30c30c",
   10293 => x"30c30c",
   10294 => x"30c30c",
   10295 => x"30c30c",
   10296 => x"30c30c",
   10297 => x"30c30c",
   10298 => x"30c30c",
   10299 => x"30c30c",
   10300 => x"30c30c",
   10301 => x"30c30c",
   10302 => x"30c30c",
   10303 => x"30c30c",
   10304 => x"30c30c",
   10305 => x"30c30c",
   10306 => x"bbffff",
   10307 => x"ffffff",
   10308 => x"ffffff",
   10309 => x"ffffff",
   10310 => x"ffffff",
   10311 => x"ffffff",
   10312 => x"ffffff",
   10313 => x"ffffff",
   10314 => x"ffffff",
   10315 => x"ffffff",
   10316 => x"ffffff",
   10317 => x"ffffff",
   10318 => x"ffffff",
   10319 => x"ffffff",
   10320 => x"ffffff",
   10321 => x"ffffff",
   10322 => x"ffffff",
   10323 => x"ffffff",
   10324 => x"ffffff",
   10325 => x"ffffff",
   10326 => x"ffffff",
   10327 => x"ffffff",
   10328 => x"ffffff",
   10329 => x"ffffff",
   10330 => x"ffffff",
   10331 => x"ffffff",
   10332 => x"ffffff",
   10333 => x"ffffff",
   10334 => x"ffffff",
   10335 => x"fffa95",
   10336 => x"abffff",
   10337 => x"ffffff",
   10338 => x"ffffff",
   10339 => x"ffffff",
   10340 => x"ffffff",
   10341 => x"ffffff",
   10342 => x"ffffff",
   10343 => x"ffffff",
   10344 => x"ffffff",
   10345 => x"ffffff",
   10346 => x"ffffff",
   10347 => x"ffffff",
   10348 => x"ffffff",
   10349 => x"ffffff",
   10350 => x"ffffff",
   10351 => x"ffffff",
   10352 => x"ffffff",
   10353 => x"ffffff",
   10354 => x"ffffff",
   10355 => x"ffffff",
   10356 => x"ffffff",
   10357 => x"ffffff",
   10358 => x"ffffff",
   10359 => x"ffffff",
   10360 => x"ffffff",
   10361 => x"ffffff",
   10362 => x"ffffff",
   10363 => x"ffffff",
   10364 => x"ffffff",
   10365 => x"ffffff",
   10366 => x"ffffff",
   10367 => x"ffffff",
   10368 => x"ffffff",
   10369 => x"ffffff",
   10370 => x"ffffff",
   10371 => x"ffffff",
   10372 => x"ffffff",
   10373 => x"ffffff",
   10374 => x"ffffff",
   10375 => x"ffffff",
   10376 => x"ffffff",
   10377 => x"ffffff",
   10378 => x"ffffff",
   10379 => x"ffffff",
   10380 => x"ffffff",
   10381 => x"ffffff",
   10382 => x"ffffff",
   10383 => x"ffffff",
   10384 => x"ffffff",
   10385 => x"ffffff",
   10386 => x"ffffff",
   10387 => x"ffffff",
   10388 => x"ffffff",
   10389 => x"ffffff",
   10390 => x"ffffff",
   10391 => x"ffffff",
   10392 => x"ffffff",
   10393 => x"ffffff",
   10394 => x"ffffff",
   10395 => x"ffffff",
   10396 => x"ffffff",
   10397 => x"ffffff",
   10398 => x"ffffff",
   10399 => x"ffffff",
   10400 => x"ffffff",
   10401 => x"ffffff",
   10402 => x"ffad70",
   10403 => x"c30c30",
   10404 => x"c30c30",
   10405 => x"c30c30",
   10406 => x"c30c30",
   10407 => x"c30c30",
   10408 => x"c30c30",
   10409 => x"c30c30",
   10410 => x"c30c30",
   10411 => x"c30c30",
   10412 => x"c30c30",
   10413 => x"c30c30",
   10414 => x"c30c30",
   10415 => x"c30c30",
   10416 => x"c30c30",
   10417 => x"c30c30",
   10418 => x"c30c30",
   10419 => x"c30c30",
   10420 => x"c30c30",
   10421 => x"c30c30",
   10422 => x"c30c30",
   10423 => x"c30c30",
   10424 => x"c28f3c",
   10425 => x"f3cf3c",
   10426 => x"f3cf3c",
   10427 => x"f3cf3c",
   10428 => x"f3cf3c",
   10429 => x"f3cf3c",
   10430 => x"f3cf3c",
   10431 => x"f3cf3c",
   10432 => x"f3cf3c",
   10433 => x"f3cf3c",
   10434 => x"f3cf3c",
   10435 => x"f3cf3c",
   10436 => x"f3cf3c",
   10437 => x"f3cf3c",
   10438 => x"f3cf3c",
   10439 => x"f3cf3c",
   10440 => x"f3cf3c",
   10441 => x"f3cf3c",
   10442 => x"f3cf3c",
   10443 => x"f3cf3c",
   10444 => x"b0c30c",
   10445 => x"30c30c",
   10446 => x"30c30c",
   10447 => x"30c30c",
   10448 => x"30c30c",
   10449 => x"30c30c",
   10450 => x"30c30c",
   10451 => x"30c30c",
   10452 => x"30c30c",
   10453 => x"30c30c",
   10454 => x"30c30c",
   10455 => x"30c30c",
   10456 => x"30c30c",
   10457 => x"30c30c",
   10458 => x"30c30c",
   10459 => x"30c30c",
   10460 => x"30c30c",
   10461 => x"30c30c",
   10462 => x"30c30c",
   10463 => x"30c30c",
   10464 => x"30c30c",
   10465 => x"30c30c",
   10466 => x"77ffff",
   10467 => x"ffffff",
   10468 => x"ffffff",
   10469 => x"ffffff",
   10470 => x"ffffff",
   10471 => x"ffffff",
   10472 => x"ffffff",
   10473 => x"ffffff",
   10474 => x"ffffff",
   10475 => x"ffffff",
   10476 => x"ffffff",
   10477 => x"ffffff",
   10478 => x"ffffff",
   10479 => x"ffffff",
   10480 => x"ffffff",
   10481 => x"ffffff",
   10482 => x"ffffff",
   10483 => x"ffffff",
   10484 => x"ffffff",
   10485 => x"ffffff",
   10486 => x"ffffff",
   10487 => x"ffffff",
   10488 => x"ffffff",
   10489 => x"ffffff",
   10490 => x"ffffff",
   10491 => x"ffffff",
   10492 => x"ffffff",
   10493 => x"ffffff",
   10494 => x"ffffff",
   10495 => x"fea56a",
   10496 => x"ffffff",
   10497 => x"ffffff",
   10498 => x"ffffff",
   10499 => x"ffffff",
   10500 => x"ffffff",
   10501 => x"ffffff",
   10502 => x"ffffff",
   10503 => x"ffffff",
   10504 => x"ffffff",
   10505 => x"ffffff",
   10506 => x"ffffff",
   10507 => x"ffffff",
   10508 => x"ffffff",
   10509 => x"ffffff",
   10510 => x"ffffff",
   10511 => x"ffffff",
   10512 => x"ffffff",
   10513 => x"ffffff",
   10514 => x"ffffff",
   10515 => x"ffffff",
   10516 => x"ffffff",
   10517 => x"ffffff",
   10518 => x"ffffff",
   10519 => x"ffffff",
   10520 => x"ffffff",
   10521 => x"ffffff",
   10522 => x"ffffff",
   10523 => x"ffffff",
   10524 => x"ffffff",
   10525 => x"ffffff",
   10526 => x"ffffff",
   10527 => x"ffffff",
   10528 => x"ffffff",
   10529 => x"ffffff",
   10530 => x"ffffff",
   10531 => x"ffffff",
   10532 => x"ffffff",
   10533 => x"ffffff",
   10534 => x"ffffff",
   10535 => x"ffffff",
   10536 => x"ffffff",
   10537 => x"ffffff",
   10538 => x"ffffff",
   10539 => x"ffffff",
   10540 => x"ffffff",
   10541 => x"ffffff",
   10542 => x"ffffff",
   10543 => x"ffffff",
   10544 => x"ffffff",
   10545 => x"ffffff",
   10546 => x"ffffff",
   10547 => x"ffffff",
   10548 => x"ffffff",
   10549 => x"ffffff",
   10550 => x"ffffff",
   10551 => x"ffffff",
   10552 => x"ffffff",
   10553 => x"ffffff",
   10554 => x"ffffff",
   10555 => x"ffffff",
   10556 => x"ffffff",
   10557 => x"ffffff",
   10558 => x"ffffff",
   10559 => x"ffffff",
   10560 => x"ffffff",
   10561 => x"ffffff",
   10562 => x"ff5c30",
   10563 => x"c30c30",
   10564 => x"c30c30",
   10565 => x"c30c30",
   10566 => x"c30c30",
   10567 => x"c30c30",
   10568 => x"c30c30",
   10569 => x"c30c30",
   10570 => x"c30c30",
   10571 => x"c30c30",
   10572 => x"c30c30",
   10573 => x"c30c30",
   10574 => x"c30c30",
   10575 => x"c30c30",
   10576 => x"c30c30",
   10577 => x"c30c30",
   10578 => x"c30c30",
   10579 => x"c30c30",
   10580 => x"c30c30",
   10581 => x"c30c30",
   10582 => x"c30c30",
   10583 => x"c30c30",
   10584 => x"92cf3c",
   10585 => x"f3cf3c",
   10586 => x"f3cf3c",
   10587 => x"f3cf3c",
   10588 => x"f3cf3c",
   10589 => x"f3cf3c",
   10590 => x"f3cf3c",
   10591 => x"f3cf3c",
   10592 => x"f3cf3c",
   10593 => x"f3cf3c",
   10594 => x"f3cf3c",
   10595 => x"f3cf3c",
   10596 => x"f3cf3c",
   10597 => x"f3cf3c",
   10598 => x"f3cf3c",
   10599 => x"f3cf3c",
   10600 => x"f3cf3c",
   10601 => x"f3cf3c",
   10602 => x"f3cf3c",
   10603 => x"f3cf3c",
   10604 => x"b1c30c",
   10605 => x"30c30c",
   10606 => x"30c30c",
   10607 => x"30c30c",
   10608 => x"30c30c",
   10609 => x"30c30c",
   10610 => x"30c30c",
   10611 => x"30c30c",
   10612 => x"30c30c",
   10613 => x"30c30c",
   10614 => x"30c30c",
   10615 => x"30c30c",
   10616 => x"30c30c",
   10617 => x"30c30c",
   10618 => x"30c30c",
   10619 => x"30c30c",
   10620 => x"30c30c",
   10621 => x"30c30c",
   10622 => x"30c30c",
   10623 => x"30c30c",
   10624 => x"30c30c",
   10625 => x"30c30c",
   10626 => x"32efff",
   10627 => x"ffffff",
   10628 => x"ffffff",
   10629 => x"ffffff",
   10630 => x"ffffff",
   10631 => x"ffffff",
   10632 => x"ffffff",
   10633 => x"ffffff",
   10634 => x"ffffff",
   10635 => x"ffffff",
   10636 => x"ffffff",
   10637 => x"ffffff",
   10638 => x"ffffff",
   10639 => x"ffffff",
   10640 => x"ffffff",
   10641 => x"ffffff",
   10642 => x"ffffff",
   10643 => x"ffffff",
   10644 => x"ffffff",
   10645 => x"ffffff",
   10646 => x"ffffff",
   10647 => x"ffffff",
   10648 => x"ffffff",
   10649 => x"ffffff",
   10650 => x"ffffff",
   10651 => x"ffffff",
   10652 => x"ffffff",
   10653 => x"ffffff",
   10654 => x"ffffff",
   10655 => x"a95abf",
   10656 => x"ffffff",
   10657 => x"ffffff",
   10658 => x"ffffff",
   10659 => x"ffffff",
   10660 => x"ffffff",
   10661 => x"ffffff",
   10662 => x"ffffff",
   10663 => x"ffffff",
   10664 => x"ffffff",
   10665 => x"ffffff",
   10666 => x"ffffff",
   10667 => x"ffffff",
   10668 => x"ffffff",
   10669 => x"ffffff",
   10670 => x"ffffff",
   10671 => x"ffffff",
   10672 => x"ffffff",
   10673 => x"ffffff",
   10674 => x"ffffff",
   10675 => x"ffffff",
   10676 => x"ffffff",
   10677 => x"ffffff",
   10678 => x"ffffff",
   10679 => x"ffffff",
   10680 => x"ffffff",
   10681 => x"ffffff",
   10682 => x"ffffff",
   10683 => x"ffffff",
   10684 => x"ffffff",
   10685 => x"ffffff",
   10686 => x"ffffff",
   10687 => x"ffffff",
   10688 => x"ffffff",
   10689 => x"ffffff",
   10690 => x"ffffff",
   10691 => x"ffffff",
   10692 => x"ffffff",
   10693 => x"ffffff",
   10694 => x"ffffff",
   10695 => x"ffffff",
   10696 => x"ffffff",
   10697 => x"ffffff",
   10698 => x"ffffff",
   10699 => x"ffffff",
   10700 => x"ffffff",
   10701 => x"ffffff",
   10702 => x"ffffff",
   10703 => x"ffffff",
   10704 => x"ffffff",
   10705 => x"ffffff",
   10706 => x"ffffff",
   10707 => x"ffffff",
   10708 => x"ffffff",
   10709 => x"ffffff",
   10710 => x"ffffff",
   10711 => x"ffffff",
   10712 => x"ffffff",
   10713 => x"ffffff",
   10714 => x"ffffff",
   10715 => x"ffffff",
   10716 => x"ffffff",
   10717 => x"ffffff",
   10718 => x"ffffff",
   10719 => x"ffffff",
   10720 => x"ffffff",
   10721 => x"ffffff",
   10722 => x"eb5c30",
   10723 => x"c30c30",
   10724 => x"c30c30",
   10725 => x"c30c30",
   10726 => x"c30c30",
   10727 => x"c30c30",
   10728 => x"c30c30",
   10729 => x"c30c30",
   10730 => x"c30c30",
   10731 => x"c30c30",
   10732 => x"c30c30",
   10733 => x"c30c30",
   10734 => x"c30c30",
   10735 => x"c30c30",
   10736 => x"c30c30",
   10737 => x"c30c30",
   10738 => x"c30c30",
   10739 => x"c30c30",
   10740 => x"c30c30",
   10741 => x"c30c30",
   10742 => x"c30c30",
   10743 => x"c30c30",
   10744 => x"a2cf3c",
   10745 => x"f3cf3c",
   10746 => x"f3cf3c",
   10747 => x"f3cf3c",
   10748 => x"f3cf3c",
   10749 => x"f3cf3c",
   10750 => x"f3cf3c",
   10751 => x"f3cf3c",
   10752 => x"f3cf3c",
   10753 => x"f3cf3c",
   10754 => x"f3cf3c",
   10755 => x"f3cf3c",
   10756 => x"f3cf3c",
   10757 => x"f3cf3c",
   10758 => x"f3cf3c",
   10759 => x"f3cf3c",
   10760 => x"f3cf3c",
   10761 => x"f3cf3c",
   10762 => x"f3cf3c",
   10763 => x"f3cf3c",
   10764 => x"f2c30c",
   10765 => x"30c30c",
   10766 => x"30c30c",
   10767 => x"30c30c",
   10768 => x"30c30c",
   10769 => x"30c30c",
   10770 => x"30c30c",
   10771 => x"30c30c",
   10772 => x"30c30c",
   10773 => x"30c30c",
   10774 => x"30c30c",
   10775 => x"30c30c",
   10776 => x"30c30c",
   10777 => x"30c30c",
   10778 => x"30c30c",
   10779 => x"30c30c",
   10780 => x"30c30c",
   10781 => x"30c30c",
   10782 => x"30c30c",
   10783 => x"30c30c",
   10784 => x"30c30c",
   10785 => x"30c30c",
   10786 => x"31dfff",
   10787 => x"ffffff",
   10788 => x"ffffff",
   10789 => x"ffffff",
   10790 => x"ffffff",
   10791 => x"ffffff",
   10792 => x"ffffff",
   10793 => x"ffffff",
   10794 => x"ffffff",
   10795 => x"ffffff",
   10796 => x"ffffff",
   10797 => x"ffffff",
   10798 => x"ffffff",
   10799 => x"ffffff",
   10800 => x"ffffff",
   10801 => x"ffffff",
   10802 => x"ffffff",
   10803 => x"ffffff",
   10804 => x"ffffff",
   10805 => x"ffffff",
   10806 => x"ffffff",
   10807 => x"ffffff",
   10808 => x"ffffff",
   10809 => x"ffffff",
   10810 => x"ffffff",
   10811 => x"ffffff",
   10812 => x"ffffff",
   10813 => x"ffffff",
   10814 => x"ffffea",
   10815 => x"56afff",
   10816 => x"ffffff",
   10817 => x"ffffff",
   10818 => x"ffffff",
   10819 => x"ffffff",
   10820 => x"ffffff",
   10821 => x"ffffff",
   10822 => x"ffffff",
   10823 => x"ffffff",
   10824 => x"ffffff",
   10825 => x"ffffff",
   10826 => x"ffffff",
   10827 => x"ffffff",
   10828 => x"ffffff",
   10829 => x"ffffff",
   10830 => x"ffffff",
   10831 => x"ffffff",
   10832 => x"ffffff",
   10833 => x"ffffff",
   10834 => x"ffffff",
   10835 => x"ffffff",
   10836 => x"ffffff",
   10837 => x"ffffff",
   10838 => x"ffffff",
   10839 => x"ffffff",
   10840 => x"ffffff",
   10841 => x"ffffff",
   10842 => x"ffffff",
   10843 => x"ffffff",
   10844 => x"ffffff",
   10845 => x"ffffff",
   10846 => x"ffffff",
   10847 => x"ffffff",
   10848 => x"ffffff",
   10849 => x"ffffff",
   10850 => x"ffffff",
   10851 => x"ffffff",
   10852 => x"ffffff",
   10853 => x"ffffff",
   10854 => x"ffffff",
   10855 => x"ffffff",
   10856 => x"ffffff",
   10857 => x"ffffff",
   10858 => x"ffffff",
   10859 => x"ffffff",
   10860 => x"ffffff",
   10861 => x"ffffff",
   10862 => x"ffffff",
   10863 => x"ffffff",
   10864 => x"ffffff",
   10865 => x"ffffff",
   10866 => x"ffffff",
   10867 => x"ffffff",
   10868 => x"ffffff",
   10869 => x"ffffff",
   10870 => x"ffffff",
   10871 => x"ffffff",
   10872 => x"ffffff",
   10873 => x"ffffff",
   10874 => x"ffffff",
   10875 => x"ffffff",
   10876 => x"ffffff",
   10877 => x"ffffff",
   10878 => x"ffffff",
   10879 => x"ffffff",
   10880 => x"ffffff",
   10881 => x"ffffff",
   10882 => x"eb0c30",
   10883 => x"c30c30",
   10884 => x"c30c30",
   10885 => x"c30c30",
   10886 => x"c30c30",
   10887 => x"c30c30",
   10888 => x"c30c30",
   10889 => x"c30c30",
   10890 => x"c30c30",
   10891 => x"c30c30",
   10892 => x"c30c30",
   10893 => x"c30c30",
   10894 => x"c30c30",
   10895 => x"c30c30",
   10896 => x"c30c30",
   10897 => x"c30c30",
   10898 => x"c30c30",
   10899 => x"c30c30",
   10900 => x"c30c30",
   10901 => x"c30c30",
   10902 => x"c30c30",
   10903 => x"c30c24",
   10904 => x"b3cf3c",
   10905 => x"f3cf3c",
   10906 => x"f3cf3c",
   10907 => x"f3cf3c",
   10908 => x"f3cf3c",
   10909 => x"f3cf3c",
   10910 => x"f3cf3c",
   10911 => x"f3cf3c",
   10912 => x"f3cf3c",
   10913 => x"f3cf3c",
   10914 => x"f3cf3c",
   10915 => x"f3cf3c",
   10916 => x"f3cf3c",
   10917 => x"f3cf3c",
   10918 => x"f3cf3c",
   10919 => x"f3cf3c",
   10920 => x"f3cf3c",
   10921 => x"f3cf3c",
   10922 => x"f3cf3c",
   10923 => x"f3cf3c",
   10924 => x"f2c70c",
   10925 => x"30c30c",
   10926 => x"30c30c",
   10927 => x"30c30c",
   10928 => x"30c30c",
   10929 => x"30c30c",
   10930 => x"30c30c",
   10931 => x"30c30c",
   10932 => x"30c30c",
   10933 => x"30c30c",
   10934 => x"30c30c",
   10935 => x"30c30c",
   10936 => x"30c30c",
   10937 => x"30c30c",
   10938 => x"30c30c",
   10939 => x"30c30c",
   10940 => x"30c30c",
   10941 => x"30c30c",
   10942 => x"30c30c",
   10943 => x"30c30c",
   10944 => x"30c30c",
   10945 => x"30c30c",
   10946 => x"30cfff",
   10947 => x"ffffff",
   10948 => x"ffffff",
   10949 => x"ffffff",
   10950 => x"ffffff",
   10951 => x"ffffff",
   10952 => x"ffffff",
   10953 => x"ffffff",
   10954 => x"ffffff",
   10955 => x"ffffff",
   10956 => x"ffffff",
   10957 => x"ffffff",
   10958 => x"ffffff",
   10959 => x"ffffff",
   10960 => x"ffffff",
   10961 => x"ffffff",
   10962 => x"ffffff",
   10963 => x"ffffff",
   10964 => x"ffffff",
   10965 => x"ffffff",
   10966 => x"ffffff",
   10967 => x"ffffff",
   10968 => x"ffffff",
   10969 => x"ffffff",
   10970 => x"ffffff",
   10971 => x"ffffff",
   10972 => x"ffffff",
   10973 => x"ffffff",
   10974 => x"fffa95",
   10975 => x"abffff",
   10976 => x"ffffff",
   10977 => x"ffffff",
   10978 => x"ffffff",
   10979 => x"ffffff",
   10980 => x"ffffff",
   10981 => x"ffffff",
   10982 => x"ffffff",
   10983 => x"ffffff",
   10984 => x"ffffff",
   10985 => x"ffffff",
   10986 => x"ffffff",
   10987 => x"ffffff",
   10988 => x"ffffff",
   10989 => x"ffffff",
   10990 => x"ffffff",
   10991 => x"ffffff",
   10992 => x"ffffff",
   10993 => x"ffffff",
   10994 => x"ffffff",
   10995 => x"ffffff",
   10996 => x"ffffff",
   10997 => x"ffffff",
   10998 => x"ffffff",
   10999 => x"ffffff",
   11000 => x"ffffff",
   11001 => x"ffffff",
   11002 => x"ffffff",
   11003 => x"ffffff",
   11004 => x"ffffff",
   11005 => x"ffffff",
   11006 => x"ffffff",
   11007 => x"ffffff",
   11008 => x"ffffff",
   11009 => x"ffffff",
   11010 => x"ffffff",
   11011 => x"ffffff",
   11012 => x"ffffff",
   11013 => x"ffffff",
   11014 => x"ffffff",
   11015 => x"ffffff",
   11016 => x"ffffff",
   11017 => x"ffffff",
   11018 => x"ffffff",
   11019 => x"ffffff",
   11020 => x"ffffff",
   11021 => x"ffffff",
   11022 => x"ffffff",
   11023 => x"ffffff",
   11024 => x"ffffff",
   11025 => x"ffffff",
   11026 => x"ffffff",
   11027 => x"ffffff",
   11028 => x"ffffff",
   11029 => x"ffffff",
   11030 => x"ffffff",
   11031 => x"ffffff",
   11032 => x"ffffff",
   11033 => x"ffffff",
   11034 => x"ffffff",
   11035 => x"ffffff",
   11036 => x"ffffff",
   11037 => x"ffffff",
   11038 => x"ffffff",
   11039 => x"ffffff",
   11040 => x"ffffff",
   11041 => x"ffffff",
   11042 => x"d70c30",
   11043 => x"c30c30",
   11044 => x"c30c30",
   11045 => x"c30c30",
   11046 => x"c30c30",
   11047 => x"c30c30",
   11048 => x"c30c30",
   11049 => x"c30c30",
   11050 => x"c30c30",
   11051 => x"c30c30",
   11052 => x"c30c30",
   11053 => x"c30c30",
   11054 => x"c30c30",
   11055 => x"c30c30",
   11056 => x"c30c30",
   11057 => x"c30c30",
   11058 => x"c30c30",
   11059 => x"c30c30",
   11060 => x"c30c30",
   11061 => x"c30c30",
   11062 => x"c30c30",
   11063 => x"c30c28",
   11064 => x"b3cf3c",
   11065 => x"f3cf3c",
   11066 => x"f3cf3c",
   11067 => x"f3cf3c",
   11068 => x"f3cf3c",
   11069 => x"f3cf3c",
   11070 => x"f3cf3c",
   11071 => x"f3cf3c",
   11072 => x"f3cf3c",
   11073 => x"f3cf3c",
   11074 => x"f3cf3c",
   11075 => x"f3cf3c",
   11076 => x"f3cf3c",
   11077 => x"f3cf3c",
   11078 => x"f3cf3c",
   11079 => x"f3cf3c",
   11080 => x"f3cf3c",
   11081 => x"f3cf3c",
   11082 => x"f3cf3c",
   11083 => x"f3cf3c",
   11084 => x"f3cb0c",
   11085 => x"30c30c",
   11086 => x"30c30c",
   11087 => x"30c30c",
   11088 => x"30c30c",
   11089 => x"30c30c",
   11090 => x"30c30c",
   11091 => x"30c30c",
   11092 => x"30c30c",
   11093 => x"30c30c",
   11094 => x"30c30c",
   11095 => x"30c30c",
   11096 => x"30c30c",
   11097 => x"30c30c",
   11098 => x"30c30c",
   11099 => x"30c30c",
   11100 => x"30c30c",
   11101 => x"30c30c",
   11102 => x"30c30c",
   11103 => x"30c30c",
   11104 => x"30c30c",
   11105 => x"30c30c",
   11106 => x"30cbbf",
   11107 => x"ffffff",
   11108 => x"ffffff",
   11109 => x"ffffff",
   11110 => x"ffffff",
   11111 => x"ffffff",
   11112 => x"ffffff",
   11113 => x"ffffff",
   11114 => x"ffffff",
   11115 => x"ffffff",
   11116 => x"ffffff",
   11117 => x"ffffff",
   11118 => x"ffffff",
   11119 => x"ffffff",
   11120 => x"ffffff",
   11121 => x"ffffff",
   11122 => x"ffffff",
   11123 => x"ffffff",
   11124 => x"ffffff",
   11125 => x"ffffff",
   11126 => x"ffffff",
   11127 => x"ffffff",
   11128 => x"ffffff",
   11129 => x"ffffff",
   11130 => x"ffffff",
   11131 => x"ffffff",
   11132 => x"ffffff",
   11133 => x"ffffff",
   11134 => x"fea56a",
   11135 => x"ffffff",
   11136 => x"ffffff",
   11137 => x"ffffff",
   11138 => x"ffffff",
   11139 => x"ffffff",
   11140 => x"ffffff",
   11141 => x"ffffff",
   11142 => x"ffffff",
   11143 => x"ffffff",
   11144 => x"ffffff",
   11145 => x"ffffff",
   11146 => x"ffffff",
   11147 => x"ffffff",
   11148 => x"ffffff",
   11149 => x"ffffff",
   11150 => x"ffffff",
   11151 => x"ffffff",
   11152 => x"ffffff",
   11153 => x"ffffff",
   11154 => x"ffffff",
   11155 => x"ffffff",
   11156 => x"ffffff",
   11157 => x"ffffff",
   11158 => x"ffffff",
   11159 => x"ffffff",
   11160 => x"ffffff",
   11161 => x"ffffff",
   11162 => x"ffffff",
   11163 => x"ffffff",
   11164 => x"ffffff",
   11165 => x"ffffff",
   11166 => x"ffffff",
   11167 => x"ffffff",
   11168 => x"ffffff",
   11169 => x"ffffff",
   11170 => x"ffffff",
   11171 => x"ffffff",
   11172 => x"ffffff",
   11173 => x"ffffff",
   11174 => x"ffffff",
   11175 => x"ffffff",
   11176 => x"ffffff",
   11177 => x"ffffff",
   11178 => x"ffffff",
   11179 => x"ffffff",
   11180 => x"ffffff",
   11181 => x"ffffff",
   11182 => x"ffffff",
   11183 => x"ffffff",
   11184 => x"ffffff",
   11185 => x"ffffff",
   11186 => x"ffffff",
   11187 => x"ffffff",
   11188 => x"ffffff",
   11189 => x"ffffff",
   11190 => x"ffffff",
   11191 => x"ffffff",
   11192 => x"ffffff",
   11193 => x"ffffff",
   11194 => x"ffffff",
   11195 => x"ffffff",
   11196 => x"ffffff",
   11197 => x"ffffff",
   11198 => x"ffffff",
   11199 => x"ffffff",
   11200 => x"ffffff",
   11201 => x"fffffa",
   11202 => x"c30c30",
   11203 => x"c30c30",
   11204 => x"c30c30",
   11205 => x"c30c30",
   11206 => x"c30c30",
   11207 => x"c30c30",
   11208 => x"c30c30",
   11209 => x"c30c30",
   11210 => x"c30c30",
   11211 => x"c30c30",
   11212 => x"c30c30",
   11213 => x"c30c30",
   11214 => x"c30c30",
   11215 => x"c30c30",
   11216 => x"c30c30",
   11217 => x"c30c30",
   11218 => x"c30c30",
   11219 => x"c30c30",
   11220 => x"c30c30",
   11221 => x"c30c30",
   11222 => x"c30c30",
   11223 => x"c30928",
   11224 => x"f3cf3c",
   11225 => x"f3cf3c",
   11226 => x"f3cf3c",
   11227 => x"f3cf3c",
   11228 => x"f3cf3c",
   11229 => x"f3cf3c",
   11230 => x"f3cf3c",
   11231 => x"f3cf3c",
   11232 => x"f3cf3c",
   11233 => x"f3cf3c",
   11234 => x"f3cf3c",
   11235 => x"f3cf3c",
   11236 => x"f3cf3c",
   11237 => x"f3cf3c",
   11238 => x"f3cf3c",
   11239 => x"f3cf3c",
   11240 => x"f3cf3c",
   11241 => x"f3cf3c",
   11242 => x"f3cf3c",
   11243 => x"f3cf3c",
   11244 => x"f3cb0c",
   11245 => x"30c30c",
   11246 => x"30c30c",
   11247 => x"30c30c",
   11248 => x"30c30c",
   11249 => x"30c30c",
   11250 => x"30c30c",
   11251 => x"30c30c",
   11252 => x"30c30c",
   11253 => x"30c30c",
   11254 => x"30c30c",
   11255 => x"30c30c",
   11256 => x"30c30c",
   11257 => x"30c30c",
   11258 => x"30c30c",
   11259 => x"30c30c",
   11260 => x"30c30c",
   11261 => x"30c30c",
   11262 => x"30c30c",
   11263 => x"30c30c",
   11264 => x"30c30c",
   11265 => x"30c30c",
   11266 => x"30c77f",
   11267 => x"ffffff",
   11268 => x"ffffff",
   11269 => x"ffffff",
   11270 => x"ffffff",
   11271 => x"ffffff",
   11272 => x"ffffff",
   11273 => x"ffffff",
   11274 => x"ffffff",
   11275 => x"ffffff",
   11276 => x"ffffff",
   11277 => x"ffffff",
   11278 => x"ffffff",
   11279 => x"ffffff",
   11280 => x"ffffff",
   11281 => x"ffffff",
   11282 => x"ffffff",
   11283 => x"ffffff",
   11284 => x"ffffff",
   11285 => x"ffffff",
   11286 => x"ffffff",
   11287 => x"ffffff",
   11288 => x"ffffff",
   11289 => x"ffffff",
   11290 => x"ffffff",
   11291 => x"ffffff",
   11292 => x"ffffff",
   11293 => x"ffffff",
   11294 => x"a95abf",
   11295 => x"ffffff",
   11296 => x"ffffff",
   11297 => x"ffffff",
   11298 => x"ffffff",
   11299 => x"ffffff",
   11300 => x"ffffff",
   11301 => x"ffffff",
   11302 => x"ffffff",
   11303 => x"ffffff",
   11304 => x"ffffff",
   11305 => x"ffffff",
   11306 => x"ffffff",
   11307 => x"ffffff",
   11308 => x"ffffff",
   11309 => x"ffffff",
   11310 => x"ffffff",
   11311 => x"ffffff",
   11312 => x"ffffff",
   11313 => x"ffffff",
   11314 => x"ffffff",
   11315 => x"ffffff",
   11316 => x"ffffff",
   11317 => x"ffffff",
   11318 => x"ffffff",
   11319 => x"ffffff",
   11320 => x"ffffff",
   11321 => x"ffffff",
   11322 => x"ffffff",
   11323 => x"ffffff",
   11324 => x"ffffff",
   11325 => x"ffffff",
   11326 => x"ffffff",
   11327 => x"ffffff",
   11328 => x"ffffff",
   11329 => x"ffffff",
   11330 => x"ffffff",
   11331 => x"ffffff",
   11332 => x"ffffff",
   11333 => x"ffffff",
   11334 => x"ffffff",
   11335 => x"ffffff",
   11336 => x"ffffff",
   11337 => x"ffffff",
   11338 => x"ffffff",
   11339 => x"ffffff",
   11340 => x"ffffff",
   11341 => x"ffffff",
   11342 => x"ffffff",
   11343 => x"ffffff",
   11344 => x"ffffff",
   11345 => x"ffffff",
   11346 => x"ffffff",
   11347 => x"ffffff",
   11348 => x"ffffff",
   11349 => x"ffffff",
   11350 => x"ffffff",
   11351 => x"ffffff",
   11352 => x"ffffff",
   11353 => x"ffffff",
   11354 => x"ffffff",
   11355 => x"ffffff",
   11356 => x"ffffff",
   11357 => x"ffffff",
   11358 => x"ffffff",
   11359 => x"ffffff",
   11360 => x"ffffff",
   11361 => x"fffff5",
   11362 => x"c30c30",
   11363 => x"c30c30",
   11364 => x"c30c30",
   11365 => x"c30c30",
   11366 => x"c30c30",
   11367 => x"c30c30",
   11368 => x"c30c30",
   11369 => x"c30c30",
   11370 => x"c30c30",
   11371 => x"c30c30",
   11372 => x"c30c30",
   11373 => x"c30c30",
   11374 => x"c30c30",
   11375 => x"c30c30",
   11376 => x"c30c30",
   11377 => x"c30c30",
   11378 => x"c30c30",
   11379 => x"c30c30",
   11380 => x"c30c30",
   11381 => x"c30c30",
   11382 => x"c30c30",
   11383 => x"c3092c",
   11384 => x"f3cf3c",
   11385 => x"f3cf3c",
   11386 => x"f3cf3c",
   11387 => x"f3cf3c",
   11388 => x"f3cf3c",
   11389 => x"f3cf3c",
   11390 => x"f3cf3c",
   11391 => x"f3cf3c",
   11392 => x"f3cf3c",
   11393 => x"f3cf3c",
   11394 => x"f3cf3c",
   11395 => x"f3cf3c",
   11396 => x"f3cf3c",
   11397 => x"f3cf3c",
   11398 => x"f3cf3c",
   11399 => x"f3cf3c",
   11400 => x"f3cf3c",
   11401 => x"f3cf3c",
   11402 => x"f3cf3c",
   11403 => x"f3cf3c",
   11404 => x"f3cf1c",
   11405 => x"30c30c",
   11406 => x"30c30c",
   11407 => x"30c30c",
   11408 => x"30c30c",
   11409 => x"30c30c",
   11410 => x"30c30c",
   11411 => x"30c30c",
   11412 => x"30c30c",
   11413 => x"30c30c",
   11414 => x"30c30c",
   11415 => x"30c30c",
   11416 => x"30c30c",
   11417 => x"30c30c",
   11418 => x"30c30c",
   11419 => x"30c30c",
   11420 => x"30c30c",
   11421 => x"30c30c",
   11422 => x"30c30c",
   11423 => x"30c30c",
   11424 => x"30c30c",
   11425 => x"30c30c",
   11426 => x"30c32e",
   11427 => x"ffffff",
   11428 => x"ffffff",
   11429 => x"ffffff",
   11430 => x"ffffff",
   11431 => x"ffffff",
   11432 => x"ffffff",
   11433 => x"ffffff",
   11434 => x"ffffff",
   11435 => x"ffffff",
   11436 => x"ffffff",
   11437 => x"ffffff",
   11438 => x"ffffff",
   11439 => x"ffffff",
   11440 => x"ffffff",
   11441 => x"ffffff",
   11442 => x"ffffff",
   11443 => x"ffffff",
   11444 => x"ffffff",
   11445 => x"ffffff",
   11446 => x"ffffff",
   11447 => x"ffffff",
   11448 => x"ffffff",
   11449 => x"ffffff",
   11450 => x"ffffff",
   11451 => x"ffffff",
   11452 => x"ffffff",
   11453 => x"ffffea",
   11454 => x"56afff",
   11455 => x"ffffff",
   11456 => x"ffffff",
   11457 => x"ffffff",
   11458 => x"ffffff",
   11459 => x"ffffff",
   11460 => x"ffffff",
   11461 => x"ffffff",
   11462 => x"ffffff",
   11463 => x"ffffff",
   11464 => x"ffffff",
   11465 => x"ffffff",
   11466 => x"ffffff",
   11467 => x"ffffff",
   11468 => x"ffffff",
   11469 => x"ffffff",
   11470 => x"ffffff",
   11471 => x"ffffff",
   11472 => x"ffffff",
   11473 => x"ffffff",
   11474 => x"ffffff",
   11475 => x"ffffff",
   11476 => x"ffffff",
   11477 => x"ffffff",
   11478 => x"ffffff",
   11479 => x"ffffff",
   11480 => x"ffffff",
   11481 => x"ffffff",
   11482 => x"ffffff",
   11483 => x"ffffff",
   11484 => x"ffffff",
   11485 => x"ffffff",
   11486 => x"ffffff",
   11487 => x"ffffff",
   11488 => x"ffffff",
   11489 => x"ffffff",
   11490 => x"ffffff",
   11491 => x"ffffff",
   11492 => x"ffffff",
   11493 => x"ffffff",
   11494 => x"ffffff",
   11495 => x"ffffff",
   11496 => x"ffffff",
   11497 => x"ffffff",
   11498 => x"ffffff",
   11499 => x"ffffff",
   11500 => x"ffffff",
   11501 => x"ffffff",
   11502 => x"ffffff",
   11503 => x"ffffff",
   11504 => x"ffffff",
   11505 => x"ffffff",
   11506 => x"ffffff",
   11507 => x"ffffff",
   11508 => x"ffffff",
   11509 => x"ffffff",
   11510 => x"ffffff",
   11511 => x"ffffff",
   11512 => x"ffffff",
   11513 => x"ffffff",
   11514 => x"ffffff",
   11515 => x"ffffff",
   11516 => x"ffffff",
   11517 => x"ffffff",
   11518 => x"ffffff",
   11519 => x"ffffff",
   11520 => x"ffffff",
   11521 => x"fffff5",
   11522 => x"c30c30",
   11523 => x"c30c30",
   11524 => x"c30c30",
   11525 => x"c30c30",
   11526 => x"c30c30",
   11527 => x"c30c30",
   11528 => x"c30c30",
   11529 => x"c30c30",
   11530 => x"c30c30",
   11531 => x"c30c30",
   11532 => x"c30c30",
   11533 => x"c30c30",
   11534 => x"c30c30",
   11535 => x"c30c30",
   11536 => x"c30c30",
   11537 => x"c30c30",
   11538 => x"c30c30",
   11539 => x"c30c30",
   11540 => x"c30c30",
   11541 => x"c30c30",
   11542 => x"c30c30",
   11543 => x"c30a2c",
   11544 => x"f3cf3c",
   11545 => x"f3cf3c",
   11546 => x"f3cf3c",
   11547 => x"f3cf3c",
   11548 => x"f3cf3c",
   11549 => x"f3cf3c",
   11550 => x"f3cf3c",
   11551 => x"f3cf3c",
   11552 => x"f3cf3c",
   11553 => x"f3cf3c",
   11554 => x"f3cf3c",
   11555 => x"f3cf3c",
   11556 => x"f3cf3c",
   11557 => x"f3cf3c",
   11558 => x"f3cf3c",
   11559 => x"f3cf3c",
   11560 => x"f3cf3c",
   11561 => x"f3cf3c",
   11562 => x"f3cf3c",
   11563 => x"f3cf3c",
   11564 => x"f3cf2c",
   11565 => x"30c30c",
   11566 => x"30c30c",
   11567 => x"30c30c",
   11568 => x"30c30c",
   11569 => x"30c30c",
   11570 => x"30c30c",
   11571 => x"30c30c",
   11572 => x"30c30c",
   11573 => x"30c30c",
   11574 => x"30c30c",
   11575 => x"30c30c",
   11576 => x"30c30c",
   11577 => x"30c30c",
   11578 => x"30c30c",
   11579 => x"30c30c",
   11580 => x"30c30c",
   11581 => x"30c30c",
   11582 => x"30c30c",
   11583 => x"30c30c",
   11584 => x"30c30c",
   11585 => x"30c30c",
   11586 => x"30c32e",
   11587 => x"ffffff",
   11588 => x"ffffff",
   11589 => x"ffffff",
   11590 => x"ffffff",
   11591 => x"ffffff",
   11592 => x"ffffff",
   11593 => x"ffffff",
   11594 => x"ffffff",
   11595 => x"ffffff",
   11596 => x"ffffff",
   11597 => x"ffffff",
   11598 => x"ffffff",
   11599 => x"ffffff",
   11600 => x"ffffff",
   11601 => x"ffffff",
   11602 => x"ffffff",
   11603 => x"ffffff",
   11604 => x"ffffff",
   11605 => x"ffffff",
   11606 => x"ffffff",
   11607 => x"ffffff",
   11608 => x"ffffff",
   11609 => x"ffffff",
   11610 => x"ffffff",
   11611 => x"ffffff",
   11612 => x"ffffff",
   11613 => x"fffa95",
   11614 => x"abffff",
   11615 => x"ffffff",
   11616 => x"ffffff",
   11617 => x"ffffff",
   11618 => x"ffffff",
   11619 => x"ffffff",
   11620 => x"ffffff",
   11621 => x"ffffff",
   11622 => x"ffffff",
   11623 => x"ffffff",
   11624 => x"ffffff",
   11625 => x"ffffff",
   11626 => x"ffffff",
   11627 => x"ffffff",
   11628 => x"ffffff",
   11629 => x"ffffff",
   11630 => x"ffffff",
   11631 => x"ffffff",
   11632 => x"ffffff",
   11633 => x"ffffff",
   11634 => x"ffffff",
   11635 => x"ffffff",
   11636 => x"ffffff",
   11637 => x"ffffff",
   11638 => x"ffffff",
   11639 => x"ffffff",
   11640 => x"ffffff",
   11641 => x"ffffff",
   11642 => x"ffffff",
   11643 => x"ffffff",
   11644 => x"ffffff",
   11645 => x"ffffff",
   11646 => x"ffffff",
   11647 => x"ffffff",
   11648 => x"ffffff",
   11649 => x"ffffff",
   11650 => x"ffffff",
   11651 => x"ffffff",
   11652 => x"ffffff",
   11653 => x"ffffff",
   11654 => x"ffffff",
   11655 => x"ffffff",
   11656 => x"ffffff",
   11657 => x"ffffff",
   11658 => x"ffffff",
   11659 => x"ffffff",
   11660 => x"ffffff",
   11661 => x"ffffff",
   11662 => x"ffffff",
   11663 => x"ffffff",
   11664 => x"ffffff",
   11665 => x"ffffff",
   11666 => x"ffffff",
   11667 => x"ffffff",
   11668 => x"ffffff",
   11669 => x"ffffff",
   11670 => x"ffffff",
   11671 => x"ffffff",
   11672 => x"ffffff",
   11673 => x"ffffff",
   11674 => x"ffffff",
   11675 => x"ffffff",
   11676 => x"ffffff",
   11677 => x"ffffff",
   11678 => x"ffffff",
   11679 => x"ffffff",
   11680 => x"ffffff",
   11681 => x"fffeb0",
   11682 => x"c30c30",
   11683 => x"c30c30",
   11684 => x"c30c30",
   11685 => x"c30c30",
   11686 => x"c30c30",
   11687 => x"c30c30",
   11688 => x"c30c30",
   11689 => x"c30c30",
   11690 => x"c30c30",
   11691 => x"c30c30",
   11692 => x"c30c30",
   11693 => x"c30c30",
   11694 => x"c30c30",
   11695 => x"c30c30",
   11696 => x"c30c30",
   11697 => x"c30c30",
   11698 => x"c30c30",
   11699 => x"c30c30",
   11700 => x"c30c30",
   11701 => x"c30c30",
   11702 => x"c30c30",
   11703 => x"c24a3c",
   11704 => x"f3cf3c",
   11705 => x"f3cf3c",
   11706 => x"f3cf3c",
   11707 => x"f3cf3c",
   11708 => x"f3cf3c",
   11709 => x"f3cf3c",
   11710 => x"f3cf3c",
   11711 => x"f3cf3c",
   11712 => x"f3cf3c",
   11713 => x"f3cf3c",
   11714 => x"f3cf3c",
   11715 => x"f3cf3c",
   11716 => x"f3cf3c",
   11717 => x"f3cf3c",
   11718 => x"f3cf3c",
   11719 => x"f3cf3c",
   11720 => x"f3cf3c",
   11721 => x"f3cf3c",
   11722 => x"f3cf3c",
   11723 => x"f3cf3c",
   11724 => x"f3cf2c",
   11725 => x"70c30c",
   11726 => x"30c30c",
   11727 => x"30c30c",
   11728 => x"30c30c",
   11729 => x"30c30c",
   11730 => x"30c30c",
   11731 => x"30c30c",
   11732 => x"30c30c",
   11733 => x"30c30c",
   11734 => x"30c30c",
   11735 => x"30c30c",
   11736 => x"30c30c",
   11737 => x"30c30c",
   11738 => x"30c30c",
   11739 => x"30c30c",
   11740 => x"30c30c",
   11741 => x"30c30c",
   11742 => x"30c30c",
   11743 => x"30c30c",
   11744 => x"30c30c",
   11745 => x"30c30c",
   11746 => x"30c31d",
   11747 => x"ffffff",
   11748 => x"ffffff",
   11749 => x"ffffff",
   11750 => x"ffffff",
   11751 => x"ffffff",
   11752 => x"ffffff",
   11753 => x"ffffff",
   11754 => x"ffffff",
   11755 => x"ffffff",
   11756 => x"ffffff",
   11757 => x"ffffff",
   11758 => x"ffffff",
   11759 => x"ffffff",
   11760 => x"ffffff",
   11761 => x"ffffff",
   11762 => x"ffffff",
   11763 => x"ffffff",
   11764 => x"ffffff",
   11765 => x"ffffff",
   11766 => x"ffffff",
   11767 => x"ffffff",
   11768 => x"ffffff",
   11769 => x"ffffff",
   11770 => x"ffffff",
   11771 => x"ffffff",
   11772 => x"ffffff",
   11773 => x"fea56a",
   11774 => x"ffffff",
   11775 => x"ffffff",
   11776 => x"ffffff",
   11777 => x"ffffff",
   11778 => x"ffffff",
   11779 => x"ffffff",
   11780 => x"ffffff",
   11781 => x"ffffff",
   11782 => x"ffffff",
   11783 => x"ffffff",
   11784 => x"ffffff",
   11785 => x"ffffff",
   11786 => x"ffffff",
   11787 => x"ffffff",
   11788 => x"ffffff",
   11789 => x"ffffff",
   11790 => x"ffffff",
   11791 => x"ffffff",
   11792 => x"ffffff",
   11793 => x"ffffff",
   11794 => x"ffffff",
   11795 => x"ffffff",
   11796 => x"ffffff",
   11797 => x"ffffff",
   11798 => x"ffffff",
   11799 => x"ffffff",
   11800 => x"ffffff",
   11801 => x"ffffff",
   11802 => x"ffffff",
   11803 => x"ffffff",
   11804 => x"ffffff",
   11805 => x"ffffff",
   11806 => x"ffffff",
   11807 => x"ffffff",
   11808 => x"ffffff",
   11809 => x"ffffff",
   11810 => x"ffffff",
   11811 => x"ffffff",
   11812 => x"ffffff",
   11813 => x"ffffff",
   11814 => x"ffffff",
   11815 => x"ffffff",
   11816 => x"ffffff",
   11817 => x"ffffff",
   11818 => x"ffffff",
   11819 => x"ffffff",
   11820 => x"ffffff",
   11821 => x"ffffff",
   11822 => x"ffffff",
   11823 => x"ffffff",
   11824 => x"ffffff",
   11825 => x"ffffff",
   11826 => x"ffffff",
   11827 => x"ffffff",
   11828 => x"ffffff",
   11829 => x"ffffff",
   11830 => x"ffffff",
   11831 => x"ffffff",
   11832 => x"ffffff",
   11833 => x"ffffff",
   11834 => x"ffffff",
   11835 => x"ffffff",
   11836 => x"ffffff",
   11837 => x"ffffff",
   11838 => x"ffffff",
   11839 => x"ffffff",
   11840 => x"ffffff",
   11841 => x"fffd70",
   11842 => x"c30c30",
   11843 => x"c30c30",
   11844 => x"c30c30",
   11845 => x"c30c30",
   11846 => x"c30c30",
   11847 => x"c30c30",
   11848 => x"c30c30",
   11849 => x"c30c30",
   11850 => x"c30c30",
   11851 => x"c30c30",
   11852 => x"c30c30",
   11853 => x"c30c30",
   11854 => x"c30c30",
   11855 => x"c30c30",
   11856 => x"c30c30",
   11857 => x"c30c30",
   11858 => x"c30c30",
   11859 => x"c30c30",
   11860 => x"c30c30",
   11861 => x"c30c30",
   11862 => x"c30c30",
   11863 => x"c24b3c",
   11864 => x"f3cf3c",
   11865 => x"f3cf3c",
   11866 => x"f3cf3c",
   11867 => x"f3cf3c",
   11868 => x"f3cf3c",
   11869 => x"f3cf3c",
   11870 => x"f3cf3c",
   11871 => x"f3cf3c",
   11872 => x"f3cf3c",
   11873 => x"f3cf3c",
   11874 => x"f3cf3c",
   11875 => x"f3cf3c",
   11876 => x"f3cf3c",
   11877 => x"f3cf3c",
   11878 => x"f3cf3c",
   11879 => x"f3cf3c",
   11880 => x"f3cf3c",
   11881 => x"f3cf3c",
   11882 => x"f3cf3c",
   11883 => x"f3cf3c",
   11884 => x"f3cf3c",
   11885 => x"70c30c",
   11886 => x"30c30c",
   11887 => x"30c30c",
   11888 => x"30c30c",
   11889 => x"30c30c",
   11890 => x"30c30c",
   11891 => x"30c30c",
   11892 => x"30c30c",
   11893 => x"30c30c",
   11894 => x"30c30c",
   11895 => x"30c30c",
   11896 => x"30c30c",
   11897 => x"30c30c",
   11898 => x"30c30c",
   11899 => x"30c30c",
   11900 => x"30c30c",
   11901 => x"30c30c",
   11902 => x"30c30c",
   11903 => x"30c30c",
   11904 => x"30c30c",
   11905 => x"30c30c",
   11906 => x"30c30c",
   11907 => x"bbffff",
   11908 => x"ffffff",
   11909 => x"ffffff",
   11910 => x"ffffff",
   11911 => x"ffffff",
   11912 => x"ffffff",
   11913 => x"ffffff",
   11914 => x"ffffff",
   11915 => x"ffffff",
   11916 => x"ffffff",
   11917 => x"ffffff",
   11918 => x"ffffff",
   11919 => x"ffffff",
   11920 => x"ffffff",
   11921 => x"ffffff",
   11922 => x"ffffff",
   11923 => x"ffffff",
   11924 => x"ffffff",
   11925 => x"ffffff",
   11926 => x"ffffff",
   11927 => x"ffffff",
   11928 => x"ffffff",
   11929 => x"ffffff",
   11930 => x"ffffff",
   11931 => x"ffffff",
   11932 => x"ffffff",
   11933 => x"a95abf",
   11934 => x"ffffff",
   11935 => x"ffffff",
   11936 => x"ffffff",
   11937 => x"ffffff",
   11938 => x"ffffff",
   11939 => x"ffffff",
   11940 => x"ffffff",
   11941 => x"ffffff",
   11942 => x"ffffff",
   11943 => x"ffffff",
   11944 => x"ffffff",
   11945 => x"ffffff",
   11946 => x"ffffff",
   11947 => x"ffffff",
   11948 => x"ffffff",
   11949 => x"ffffff",
   11950 => x"ffffff",
   11951 => x"ffffff",
   11952 => x"ffffff",
   11953 => x"ffffff",
   11954 => x"ffffff",
   11955 => x"ffffff",
   11956 => x"ffffff",
   11957 => x"ffffff",
   11958 => x"ffffff",
   11959 => x"ffffff",
   11960 => x"ffffff",
   11961 => x"ffffff",
   11962 => x"ffffff",
   11963 => x"ffffff",
   11964 => x"ffffff",
   11965 => x"ffffff",
   11966 => x"ffffff",
   11967 => x"ffffff",
   11968 => x"ffffff",
   11969 => x"ffffff",
   11970 => x"ffffff",
   11971 => x"ffffff",
   11972 => x"ffffff",
   11973 => x"ffffff",
   11974 => x"ffffff",
   11975 => x"ffffff",
   11976 => x"ffffff",
   11977 => x"ffffff",
   11978 => x"ffffff",
   11979 => x"ffffff",
   11980 => x"ffffff",
   11981 => x"ffffff",
   11982 => x"ffffff",
   11983 => x"ffffff",
   11984 => x"ffffff",
   11985 => x"ffffff",
   11986 => x"ffffff",
   11987 => x"ffffff",
   11988 => x"ffffff",
   11989 => x"ffffff",
   11990 => x"ffffff",
   11991 => x"ffffff",
   11992 => x"ffffff",
   11993 => x"ffffff",
   11994 => x"ffffff",
   11995 => x"ffffff",
   11996 => x"ffffff",
   11997 => x"ffffff",
   11998 => x"ffffff",
   11999 => x"ffffff",
   12000 => x"ffffff",
   12001 => x"fffd70",
   12002 => x"c30c30",
   12003 => x"c30c30",
   12004 => x"c30c30",
   12005 => x"c30c30",
   12006 => x"c30c30",
   12007 => x"c30c30",
   12008 => x"c30c30",
   12009 => x"c30c30",
   12010 => x"c30c30",
   12011 => x"c30c30",
   12012 => x"c30c30",
   12013 => x"c30c30",
   12014 => x"c30c30",
   12015 => x"c30c30",
   12016 => x"c30c30",
   12017 => x"c30c30",
   12018 => x"c30c30",
   12019 => x"c30c30",
   12020 => x"c30c30",
   12021 => x"c30c30",
   12022 => x"c30c30",
   12023 => x"c28b3c",
   12024 => x"f3cf3c",
   12025 => x"f3cf3c",
   12026 => x"f3cf3c",
   12027 => x"f3cf3c",
   12028 => x"f3cf3c",
   12029 => x"f3cf3c",
   12030 => x"f3cf3c",
   12031 => x"f3cf3c",
   12032 => x"f3cf3c",
   12033 => x"f3cf3c",
   12034 => x"f3cf3c",
   12035 => x"f3cf3c",
   12036 => x"f3cf3c",
   12037 => x"f3cf3c",
   12038 => x"f3cf3c",
   12039 => x"f3cf3c",
   12040 => x"f3cf3c",
   12041 => x"f3cf3c",
   12042 => x"f3cf3c",
   12043 => x"f3cf3c",
   12044 => x"f3cf3c",
   12045 => x"b0c30c",
   12046 => x"30c30c",
   12047 => x"30c30c",
   12048 => x"30c30c",
   12049 => x"30c30c",
   12050 => x"30c30c",
   12051 => x"30c30c",
   12052 => x"30c30c",
   12053 => x"30c30c",
   12054 => x"30c30c",
   12055 => x"30c30c",
   12056 => x"30c30c",
   12057 => x"30c30c",
   12058 => x"30c30c",
   12059 => x"30c30c",
   12060 => x"30c30c",
   12061 => x"30c30c",
   12062 => x"30c30c",
   12063 => x"30c30c",
   12064 => x"30c30c",
   12065 => x"30c30c",
   12066 => x"30c30c",
   12067 => x"77ffff",
   12068 => x"ffffff",
   12069 => x"ffffff",
   12070 => x"ffffff",
   12071 => x"ffffff",
   12072 => x"ffffff",
   12073 => x"ffffff",
   12074 => x"ffffff",
   12075 => x"ffffff",
   12076 => x"ffffff",
   12077 => x"ffffff",
   12078 => x"ffffff",
   12079 => x"ffffff",
   12080 => x"ffffff",
   12081 => x"ffffff",
   12082 => x"ffffff",
   12083 => x"ffffff",
   12084 => x"ffffff",
   12085 => x"ffffff",
   12086 => x"ffffff",
   12087 => x"ffffff",
   12088 => x"ffffff",
   12089 => x"ffffff",
   12090 => x"ffffff",
   12091 => x"ffffff",
   12092 => x"ffffea",
   12093 => x"56afff",
   12094 => x"ffffff",
   12095 => x"ffffff",
   12096 => x"ffffff",
   12097 => x"ffffff",
   12098 => x"ffffff",
   12099 => x"ffffff",
   12100 => x"ffffff",
   12101 => x"ffffff",
   12102 => x"ffffff",
   12103 => x"ffffff",
   12104 => x"ffffff",
   12105 => x"ffffff",
   12106 => x"ffffff",
   12107 => x"ffffff",
   12108 => x"ffffff",
   12109 => x"ffffff",
   12110 => x"ffffff",
   12111 => x"ffffff",
   12112 => x"ffffff",
   12113 => x"ffffff",
   12114 => x"ffffff",
   12115 => x"ffffff",
   12116 => x"ffffff",
   12117 => x"ffffff",
   12118 => x"ffffff",
   12119 => x"ffffff",
   12120 => x"ffffff",
   12121 => x"ffffff",
   12122 => x"ffffff",
   12123 => x"ffffff",
   12124 => x"ffffff",
   12125 => x"ffffff",
   12126 => x"ffffff",
   12127 => x"ffffff",
   12128 => x"ffffff",
   12129 => x"ffffff",
   12130 => x"ffffff",
   12131 => x"ffffff",
   12132 => x"ffffff",
   12133 => x"ffffff",
   12134 => x"ffffff",
   12135 => x"ffffff",
   12136 => x"ffffff",
   12137 => x"ffffff",
   12138 => x"ffffff",
   12139 => x"ffffff",
   12140 => x"ffffff",
   12141 => x"ffffff",
   12142 => x"ffffff",
   12143 => x"ffffff",
   12144 => x"ffffff",
   12145 => x"ffffff",
   12146 => x"ffffff",
   12147 => x"ffffff",
   12148 => x"ffffff",
   12149 => x"ffffff",
   12150 => x"ffffff",
   12151 => x"ffffff",
   12152 => x"ffffff",
   12153 => x"ffffff",
   12154 => x"ffffff",
   12155 => x"ffffff",
   12156 => x"ffffff",
   12157 => x"ffffff",
   12158 => x"ffffff",
   12159 => x"ffffff",
   12160 => x"ffffff",
   12161 => x"ffac30",
   12162 => x"c30c30",
   12163 => x"c30c30",
   12164 => x"c30c30",
   12165 => x"c30c30",
   12166 => x"c30c30",
   12167 => x"c30c30",
   12168 => x"c30c30",
   12169 => x"c30c30",
   12170 => x"c30c30",
   12171 => x"c30c30",
   12172 => x"c30c30",
   12173 => x"c30c30",
   12174 => x"c30c30",
   12175 => x"c30c30",
   12176 => x"c30c30",
   12177 => x"c30c30",
   12178 => x"c30c30",
   12179 => x"c30c30",
   12180 => x"c30c30",
   12181 => x"c30c30",
   12182 => x"c30c30",
   12183 => x"92cf3c",
   12184 => x"f3cf3c",
   12185 => x"f3cf3c",
   12186 => x"f3cf3c",
   12187 => x"f3cf3c",
   12188 => x"f3cf3c",
   12189 => x"f3cf3c",
   12190 => x"f3cf3c",
   12191 => x"f3cf3c",
   12192 => x"f3cf3c",
   12193 => x"f3cf3c",
   12194 => x"f3cf3c",
   12195 => x"f3cf3c",
   12196 => x"f3cf3c",
   12197 => x"f3cf3c",
   12198 => x"f3cf3c",
   12199 => x"f3cf3c",
   12200 => x"f3cf3c",
   12201 => x"f3cf3c",
   12202 => x"f3cf3c",
   12203 => x"f3cf3c",
   12204 => x"f3cf3c",
   12205 => x"f1c30c",
   12206 => x"30c30c",
   12207 => x"30c30c",
   12208 => x"30c30c",
   12209 => x"30c30c",
   12210 => x"30c30c",
   12211 => x"30c30c",
   12212 => x"30c30c",
   12213 => x"30c30c",
   12214 => x"30c30c",
   12215 => x"30c30c",
   12216 => x"30c30c",
   12217 => x"30c30c",
   12218 => x"30c30c",
   12219 => x"30c30c",
   12220 => x"30c30c",
   12221 => x"30c30c",
   12222 => x"30c30c",
   12223 => x"30c30c",
   12224 => x"30c30c",
   12225 => x"30c30c",
   12226 => x"30c30c",
   12227 => x"33ffff",
   12228 => x"ffffff",
   12229 => x"ffffff",
   12230 => x"ffffff",
   12231 => x"ffffff",
   12232 => x"ffffff",
   12233 => x"ffffff",
   12234 => x"ffffff",
   12235 => x"ffffff",
   12236 => x"ffffff",
   12237 => x"ffffff",
   12238 => x"ffffff",
   12239 => x"ffffff",
   12240 => x"ffffff",
   12241 => x"ffffff",
   12242 => x"ffffff",
   12243 => x"ffffff",
   12244 => x"ffffff",
   12245 => x"ffffff",
   12246 => x"ffffff",
   12247 => x"ffffff",
   12248 => x"ffffff",
   12249 => x"ffffff",
   12250 => x"ffffff",
   12251 => x"ffffff",
   12252 => x"fffa95",
   12253 => x"abffff",
   12254 => x"ffffff",
   12255 => x"ffffff",
   12256 => x"ffffff",
   12257 => x"ffffff",
   12258 => x"ffffff",
   12259 => x"ffffff",
   12260 => x"ffffff",
   12261 => x"ffffff",
   12262 => x"ffffff",
   12263 => x"ffffff",
   12264 => x"ffffff",
   12265 => x"ffffff",
   12266 => x"ffffff",
   12267 => x"ffffff",
   12268 => x"ffffff",
   12269 => x"ffffff",
   12270 => x"ffffff",
   12271 => x"ffffff",
   12272 => x"ffffff",
   12273 => x"ffffff",
   12274 => x"ffffff",
   12275 => x"ffffff",
   12276 => x"ffffff",
   12277 => x"ffffff",
   12278 => x"ffffff",
   12279 => x"ffffff",
   12280 => x"ffffff",
   12281 => x"ffffff",
   12282 => x"ffffff",
   12283 => x"ffffff",
   12284 => x"ffffff",
   12285 => x"ffffff",
   12286 => x"ffffff",
   12287 => x"ffffff",
   12288 => x"ffffff",
   12289 => x"ffffff",
   12290 => x"ffffff",
   12291 => x"ffffff",
   12292 => x"ffffff",
   12293 => x"ffffff",
   12294 => x"ffffff",
   12295 => x"ffffff",
   12296 => x"ffffff",
   12297 => x"ffffff",
   12298 => x"ffffff",
   12299 => x"ffffff",
   12300 => x"ffffff",
   12301 => x"ffffff",
   12302 => x"ffffff",
   12303 => x"ffffff",
   12304 => x"ffffff",
   12305 => x"ffffff",
   12306 => x"ffffff",
   12307 => x"ffffff",
   12308 => x"ffffff",
   12309 => x"ffffff",
   12310 => x"ffffff",
   12311 => x"ffffff",
   12312 => x"ffffff",
   12313 => x"ffffff",
   12314 => x"ffffff",
   12315 => x"ffffff",
   12316 => x"ffffff",
   12317 => x"ffffff",
   12318 => x"ffffff",
   12319 => x"ffffff",
   12320 => x"ffffff",
   12321 => x"ff5c30",
   12322 => x"c30c30",
   12323 => x"c30c30",
   12324 => x"c30c30",
   12325 => x"c30c30",
   12326 => x"c30c30",
   12327 => x"c30c30",
   12328 => x"c30c30",
   12329 => x"c30c30",
   12330 => x"c30c30",
   12331 => x"c30c30",
   12332 => x"c30c30",
   12333 => x"c30c30",
   12334 => x"c30c30",
   12335 => x"c30c30",
   12336 => x"c30c30",
   12337 => x"c30c30",
   12338 => x"c30c30",
   12339 => x"c30c30",
   12340 => x"c30c30",
   12341 => x"c30c30",
   12342 => x"c30c30",
   12343 => x"a2cf3c",
   12344 => x"f3cf3c",
   12345 => x"f3cf3c",
   12346 => x"f3cf3c",
   12347 => x"f3cf3c",
   12348 => x"f3cf3c",
   12349 => x"f3cf3c",
   12350 => x"f3cf3c",
   12351 => x"f3cf3c",
   12352 => x"f3cf3c",
   12353 => x"f3cf3c",
   12354 => x"f3cf3c",
   12355 => x"f3cf3c",
   12356 => x"f3cf3c",
   12357 => x"f3cf3c",
   12358 => x"f3cf3c",
   12359 => x"f3cf3c",
   12360 => x"f3cf3c",
   12361 => x"f3cf3c",
   12362 => x"f3cf3c",
   12363 => x"f3cf3c",
   12364 => x"f3cf3c",
   12365 => x"f2c30c",
   12366 => x"30c30c",
   12367 => x"30c30c",
   12368 => x"30c30c",
   12369 => x"30c30c",
   12370 => x"30c30c",
   12371 => x"30c30c",
   12372 => x"30c30c",
   12373 => x"30c30c",
   12374 => x"30c30c",
   12375 => x"30c30c",
   12376 => x"30c30c",
   12377 => x"30c30c",
   12378 => x"30c30c",
   12379 => x"30c30c",
   12380 => x"30c30c",
   12381 => x"30c30c",
   12382 => x"30c30c",
   12383 => x"30c30c",
   12384 => x"30c30c",
   12385 => x"30c30c",
   12386 => x"30c30c",
   12387 => x"32efff",
   12388 => x"ffffff",
   12389 => x"ffffff",
   12390 => x"ffffff",
   12391 => x"ffffff",
   12392 => x"ffffff",
   12393 => x"ffffff",
   12394 => x"ffffff",
   12395 => x"ffffff",
   12396 => x"ffffff",
   12397 => x"ffffff",
   12398 => x"ffffff",
   12399 => x"ffffff",
   12400 => x"ffffff",
   12401 => x"ffffff",
   12402 => x"ffffff",
   12403 => x"ffffff",
   12404 => x"ffffff",
   12405 => x"ffffff",
   12406 => x"ffffff",
   12407 => x"ffffff",
   12408 => x"ffffff",
   12409 => x"ffffff",
   12410 => x"ffffff",
   12411 => x"ffffff",
   12412 => x"fea56a",
   12413 => x"ffffff",
   12414 => x"ffffff",
   12415 => x"ffffff",
   12416 => x"ffffff",
   12417 => x"ffffff",
   12418 => x"ffffff",
   12419 => x"ffffff",
   12420 => x"ffffff",
   12421 => x"ffffff",
   12422 => x"ffffff",
   12423 => x"ffffff",
   12424 => x"ffffff",
   12425 => x"ffffff",
   12426 => x"ffffff",
   12427 => x"ffffff",
   12428 => x"ffffff",
   12429 => x"ffffff",
   12430 => x"ffffff",
   12431 => x"ffffff",
   12432 => x"ffffff",
   12433 => x"ffffff",
   12434 => x"ffffff",
   12435 => x"ffffff",
   12436 => x"ffffff",
   12437 => x"ffffff",
   12438 => x"ffffff",
   12439 => x"ffffff",
   12440 => x"ffffff",
   12441 => x"ffffff",
   12442 => x"ffffff",
   12443 => x"ffffff",
   12444 => x"ffffff",
   12445 => x"ffffff",
   12446 => x"ffffff",
   12447 => x"ffffff",
   12448 => x"ffffff",
   12449 => x"ffffff",
   12450 => x"ffffff",
   12451 => x"ffffff",
   12452 => x"ffffff",
   12453 => x"ffffff",
   12454 => x"ffffff",
   12455 => x"ffffff",
   12456 => x"ffffff",
   12457 => x"ffffff",
   12458 => x"ffffff",
   12459 => x"ffffff",
   12460 => x"ffffff",
   12461 => x"ffffff",
   12462 => x"ffffff",
   12463 => x"ffffff",
   12464 => x"ffffff",
   12465 => x"ffffff",
   12466 => x"ffffff",
   12467 => x"ffffff",
   12468 => x"ffffff",
   12469 => x"ffffff",
   12470 => x"ffffff",
   12471 => x"ffffff",
   12472 => x"ffffff",
   12473 => x"ffffff",
   12474 => x"ffffff",
   12475 => x"ffffff",
   12476 => x"ffffff",
   12477 => x"ffffff",
   12478 => x"ffffff",
   12479 => x"ffffff",
   12480 => x"ffffff",
   12481 => x"ff5c30",
   12482 => x"c30c30",
   12483 => x"c30c30",
   12484 => x"c30c30",
   12485 => x"c30c30",
   12486 => x"c30c30",
   12487 => x"c30c30",
   12488 => x"c30c30",
   12489 => x"c30c30",
   12490 => x"c30c30",
   12491 => x"c30c30",
   12492 => x"c30c30",
   12493 => x"c30c30",
   12494 => x"c30c30",
   12495 => x"c30c30",
   12496 => x"c30c30",
   12497 => x"c30c30",
   12498 => x"c30c30",
   12499 => x"c30c30",
   12500 => x"c30c30",
   12501 => x"c30c30",
   12502 => x"c30c30",
   12503 => x"a2cf3c",
   12504 => x"f3cf3c",
   12505 => x"f3cf3c",
   12506 => x"f3cf3c",
   12507 => x"f3cf3c",
   12508 => x"f3cf3c",
   12509 => x"f3cf3c",
   12510 => x"f3cf3c",
   12511 => x"f3cf3c",
   12512 => x"f3cf3c",
   12513 => x"f3cf3c",
   12514 => x"f3cf3c",
   12515 => x"f3cf3c",
   12516 => x"f3cf3c",
   12517 => x"f3cf3c",
   12518 => x"f3cf3c",
   12519 => x"f3cf3c",
   12520 => x"f3cf3c",
   12521 => x"f3cf3c",
   12522 => x"f3cf3c",
   12523 => x"f3cf3c",
   12524 => x"f3cf3c",
   12525 => x"f2c30c",
   12526 => x"30c30c",
   12527 => x"30c30c",
   12528 => x"30c30c",
   12529 => x"30c30c",
   12530 => x"30c30c",
   12531 => x"30c30c",
   12532 => x"30c30c",
   12533 => x"30c30c",
   12534 => x"30c30c",
   12535 => x"30c30c",
   12536 => x"30c30c",
   12537 => x"30c30c",
   12538 => x"30c30c",
   12539 => x"30c30c",
   12540 => x"30c30c",
   12541 => x"30c30c",
   12542 => x"30c30c",
   12543 => x"30c30c",
   12544 => x"30c30c",
   12545 => x"30c30c",
   12546 => x"30c30c",
   12547 => x"31dfff",
   12548 => x"ffffff",
   12549 => x"ffffff",
   12550 => x"ffffff",
   12551 => x"ffffff",
   12552 => x"ffffff",
   12553 => x"ffffff",
   12554 => x"ffffff",
   12555 => x"ffffff",
   12556 => x"ffffff",
   12557 => x"ffffff",
   12558 => x"ffffff",
   12559 => x"ffffff",
   12560 => x"ffffff",
   12561 => x"ffffff",
   12562 => x"ffffff",
   12563 => x"ffffff",
   12564 => x"ffffff",
   12565 => x"ffffff",
   12566 => x"ffffff",
   12567 => x"ffffff",
   12568 => x"ffffff",
   12569 => x"ffffff",
   12570 => x"ffffff",
   12571 => x"ffffff",
   12572 => x"a95abf",
   12573 => x"ffffff",
   12574 => x"ffffff",
   12575 => x"ffffff",
   12576 => x"ffffff",
   12577 => x"ffffff",
   12578 => x"ffffff",
   12579 => x"ffffff",
   12580 => x"ffffff",
   12581 => x"ffffff",
   12582 => x"ffffff",
   12583 => x"ffffff",
   12584 => x"ffffff",
   12585 => x"ffffff",
   12586 => x"ffffff",
   12587 => x"ffffff",
   12588 => x"ffffff",
   12589 => x"ffffff",
   12590 => x"ffffff",
   12591 => x"ffffff",
   12592 => x"ffffff",
   12593 => x"ffffff",
   12594 => x"ffffff",
   12595 => x"ffffff",
   12596 => x"ffffff",
   12597 => x"ffffff",
   12598 => x"ffffff",
   12599 => x"ffffff",
   12600 => x"ffffff",
   12601 => x"ffffff",
   12602 => x"ffffff",
   12603 => x"ffffff",
   12604 => x"ffffff",
   12605 => x"ffffff",
   12606 => x"ffffff",
   12607 => x"ffffff",
   12608 => x"ffffff",
   12609 => x"ffffff",
   12610 => x"ffffff",
   12611 => x"ffffff",
   12612 => x"ffffff",
   12613 => x"ffffff",
   12614 => x"ffffff",
   12615 => x"ffffff",
   12616 => x"ffffff",
   12617 => x"ffffff",
   12618 => x"ffffff",
   12619 => x"ffffff",
   12620 => x"ffffff",
   12621 => x"ffffff",
   12622 => x"ffffff",
   12623 => x"ffffff",
   12624 => x"ffffff",
   12625 => x"ffffff",
   12626 => x"ffffff",
   12627 => x"ffffff",
   12628 => x"ffffff",
   12629 => x"ffffff",
   12630 => x"ffffff",
   12631 => x"ffffff",
   12632 => x"ffffff",
   12633 => x"ffffff",
   12634 => x"ffffff",
   12635 => x"ffffff",
   12636 => x"ffffff",
   12637 => x"ffffff",
   12638 => x"ffffff",
   12639 => x"ffffff",
   12640 => x"ffffff",
   12641 => x"eb0c30",
   12642 => x"c30c30",
   12643 => x"c30c30",
   12644 => x"c30c30",
   12645 => x"c30c30",
   12646 => x"c30c30",
   12647 => x"c30c30",
   12648 => x"c30c30",
   12649 => x"c30c30",
   12650 => x"c30c30",
   12651 => x"c30c30",
   12652 => x"c30c30",
   12653 => x"c30c30",
   12654 => x"c30c30",
   12655 => x"c30c30",
   12656 => x"c30c30",
   12657 => x"c30c30",
   12658 => x"c30c30",
   12659 => x"c30c30",
   12660 => x"c30c30",
   12661 => x"c30c30",
   12662 => x"c30c24",
   12663 => x"a3cf3c",
   12664 => x"f3cf3c",
   12665 => x"f3cf3c",
   12666 => x"f3cf3c",
   12667 => x"f3cf3c",
   12668 => x"f3cf3c",
   12669 => x"f3cf3c",
   12670 => x"f3cf3c",
   12671 => x"f3cf3c",
   12672 => x"f3cf3c",
   12673 => x"f3cf3c",
   12674 => x"f3cf3c",
   12675 => x"f3cf3c",
   12676 => x"f3cf3c",
   12677 => x"f3cf3c",
   12678 => x"f3cf3c",
   12679 => x"f3cf3c",
   12680 => x"f3cf3c",
   12681 => x"f3cf3c",
   12682 => x"f3cf3c",
   12683 => x"f3cf3c",
   12684 => x"f3cf3c",
   12685 => x"f3c70c",
   12686 => x"30c30c",
   12687 => x"30c30c",
   12688 => x"30c30c",
   12689 => x"30c30c",
   12690 => x"30c30c",
   12691 => x"30c30c",
   12692 => x"30c30c",
   12693 => x"30c30c",
   12694 => x"30c30c",
   12695 => x"30c30c",
   12696 => x"30c30c",
   12697 => x"30c30c",
   12698 => x"30c30c",
   12699 => x"30c30c",
   12700 => x"30c30c",
   12701 => x"30c30c",
   12702 => x"30c30c",
   12703 => x"30c30c",
   12704 => x"30c30c",
   12705 => x"30c30c",
   12706 => x"30c30c",
   12707 => x"31dfff",
   12708 => x"ffffff",
   12709 => x"ffffff",
   12710 => x"ffffff",
   12711 => x"ffffff",
   12712 => x"ffffff",
   12713 => x"ffffff",
   12714 => x"ffffff",
   12715 => x"ffffff",
   12716 => x"ffffff",
   12717 => x"ffffff",
   12718 => x"ffffff",
   12719 => x"ffffff",
   12720 => x"ffffff",
   12721 => x"ffffff",
   12722 => x"ffffff",
   12723 => x"ffffff",
   12724 => x"ffffff",
   12725 => x"ffffff",
   12726 => x"ffffff",
   12727 => x"ffffff",
   12728 => x"ffffff",
   12729 => x"ffffff",
   12730 => x"ffffff",
   12731 => x"ffffea",
   12732 => x"56afff",
   12733 => x"ffffff",
   12734 => x"ffffff",
   12735 => x"ffffff",
   12736 => x"ffffff",
   12737 => x"ffffff",
   12738 => x"ffffff",
   12739 => x"ffffff",
   12740 => x"ffffff",
   12741 => x"ffffff",
   12742 => x"ffffff",
   12743 => x"ffffff",
   12744 => x"ffffff",
   12745 => x"ffffff",
   12746 => x"ffffff",
   12747 => x"ffffff",
   12748 => x"ffffff",
   12749 => x"ffffff",
   12750 => x"ffffff",
   12751 => x"ffffff",
   12752 => x"ffffff",
   12753 => x"ffffff",
   12754 => x"ffffff",
   12755 => x"ffffff",
   12756 => x"ffffff",
   12757 => x"ffffff",
   12758 => x"ffffff",
   12759 => x"ffffff",
   12760 => x"ffffff",
   12761 => x"ffffff",
   12762 => x"ffffff",
   12763 => x"ffffff",
   12764 => x"ffffff",
   12765 => x"ffffff",
   12766 => x"ffffff",
   12767 => x"ffffff",
   12768 => x"ffffff",
   12769 => x"ffffff",
   12770 => x"ffffff",
   12771 => x"ffffff",
   12772 => x"ffffff",
   12773 => x"ffffff",
   12774 => x"ffffff",
   12775 => x"ffffff",
   12776 => x"ffffff",
   12777 => x"ffffff",
   12778 => x"ffffff",
   12779 => x"ffffff",
   12780 => x"ffffff",
   12781 => x"ffffff",
   12782 => x"ffffff",
   12783 => x"ffffff",
   12784 => x"ffffff",
   12785 => x"ffffff",
   12786 => x"ffffff",
   12787 => x"ffffff",
   12788 => x"ffffff",
   12789 => x"ffffff",
   12790 => x"ffffff",
   12791 => x"ffffff",
   12792 => x"ffffff",
   12793 => x"ffffff",
   12794 => x"ffffff",
   12795 => x"ffffff",
   12796 => x"ffffff",
   12797 => x"ffffff",
   12798 => x"ffffff",
   12799 => x"ffffff",
   12800 => x"ffffff",
   12801 => x"d70c30",
   12802 => x"c30c30",
   12803 => x"c30c30",
   12804 => x"c30c30",
   12805 => x"c30c30",
   12806 => x"c30c30",
   12807 => x"c30c30",
   12808 => x"c30c30",
   12809 => x"c30c30",
   12810 => x"c30c30",
   12811 => x"c30c30",
   12812 => x"c30c30",
   12813 => x"c30c30",
   12814 => x"c30c30",
   12815 => x"c30c30",
   12816 => x"c30c30",
   12817 => x"c30c30",
   12818 => x"c30c30",
   12819 => x"c30c30",
   12820 => x"c30c30",
   12821 => x"c30c30",
   12822 => x"c30c24",
   12823 => x"b3cf3c",
   12824 => x"f3cf3c",
   12825 => x"f3cf3c",
   12826 => x"f3cf3c",
   12827 => x"f3cf3c",
   12828 => x"f3cf3c",
   12829 => x"f3cf3c",
   12830 => x"f3cf3c",
   12831 => x"f3cf3c",
   12832 => x"f3cf3c",
   12833 => x"f3cf3c",
   12834 => x"f3cf3c",
   12835 => x"f3cf3c",
   12836 => x"f3cf3c",
   12837 => x"f3cf3c",
   12838 => x"f3cf3c",
   12839 => x"f3cf3c",
   12840 => x"f3cf3c",
   12841 => x"f3cf3c",
   12842 => x"f3cf3c",
   12843 => x"f3cf3c",
   12844 => x"f3cf3c",
   12845 => x"f3c70c",
   12846 => x"30c30c",
   12847 => x"30c30c",
   12848 => x"30c30c",
   12849 => x"30c30c",
   12850 => x"30c30c",
   12851 => x"30c30c",
   12852 => x"30c30c",
   12853 => x"30c30c",
   12854 => x"30c30c",
   12855 => x"30c30c",
   12856 => x"30c30c",
   12857 => x"30c30c",
   12858 => x"30c30c",
   12859 => x"30c30c",
   12860 => x"30c30c",
   12861 => x"30c30c",
   12862 => x"30c30c",
   12863 => x"30c30c",
   12864 => x"30c30c",
   12865 => x"30c30c",
   12866 => x"30c30c",
   12867 => x"30cfff",
   12868 => x"ffffff",
   12869 => x"ffffff",
   12870 => x"ffffff",
   12871 => x"ffffff",
   12872 => x"ffffff",
   12873 => x"ffffff",
   12874 => x"ffffff",
   12875 => x"ffffff",
   12876 => x"ffffff",
   12877 => x"ffffff",
   12878 => x"ffffff",
   12879 => x"ffffff",
   12880 => x"ffffff",
   12881 => x"ffffff",
   12882 => x"ffffff",
   12883 => x"ffffff",
   12884 => x"ffffff",
   12885 => x"ffffff",
   12886 => x"ffffff",
   12887 => x"ffffff",
   12888 => x"ffffff",
   12889 => x"ffffff",
   12890 => x"ffffff",
   12891 => x"fffa95",
   12892 => x"abffff",
   12893 => x"ffffff",
   12894 => x"ffffff",
   12895 => x"ffffff",
   12896 => x"ffffff",
   12897 => x"ffffff",
   12898 => x"ffffff",
   12899 => x"ffffff",
   12900 => x"ffffff",
   12901 => x"ffffff",
   12902 => x"ffffff",
   12903 => x"ffffff",
   12904 => x"ffffff",
   12905 => x"ffffff",
   12906 => x"ffffff",
   12907 => x"ffffff",
   12908 => x"ffffff",
   12909 => x"ffffff",
   12910 => x"ffffff",
   12911 => x"ffffff",
   12912 => x"ffffff",
   12913 => x"ffffff",
   12914 => x"ffffff",
   12915 => x"ffffff",
   12916 => x"ffffff",
   12917 => x"ffffff",
   12918 => x"ffffff",
   12919 => x"ffffff",
   12920 => x"ffffff",
   12921 => x"ffffff",
   12922 => x"ffffff",
   12923 => x"ffffff",
   12924 => x"ffffff",
   12925 => x"ffffff",
   12926 => x"ffffff",
   12927 => x"ffffff",
   12928 => x"ffffff",
   12929 => x"ffffff",
   12930 => x"ffffff",
   12931 => x"ffffff",
   12932 => x"ffffff",
   12933 => x"ffffff",
   12934 => x"ffffff",
   12935 => x"ffffff",
   12936 => x"ffffff",
   12937 => x"ffffff",
   12938 => x"ffffff",
   12939 => x"ffffff",
   12940 => x"ffffff",
   12941 => x"ffffff",
   12942 => x"ffffff",
   12943 => x"ffffff",
   12944 => x"ffffff",
   12945 => x"ffffff",
   12946 => x"ffffff",
   12947 => x"ffffff",
   12948 => x"ffffff",
   12949 => x"ffffff",
   12950 => x"ffffff",
   12951 => x"ffffff",
   12952 => x"ffffff",
   12953 => x"ffffff",
   12954 => x"ffffff",
   12955 => x"ffffff",
   12956 => x"ffffff",
   12957 => x"ffffff",
   12958 => x"ffffff",
   12959 => x"ffffff",
   12960 => x"ffffff",
   12961 => x"d70c30",
   12962 => x"c30c30",
   12963 => x"c30c30",
   12964 => x"c30c30",
   12965 => x"c30c30",
   12966 => x"c30c30",
   12967 => x"c30c30",
   12968 => x"c30c30",
   12969 => x"c30c30",
   12970 => x"c30c30",
   12971 => x"c30c30",
   12972 => x"c30c30",
   12973 => x"c30c30",
   12974 => x"c30c30",
   12975 => x"c30c30",
   12976 => x"c30c30",
   12977 => x"c30c30",
   12978 => x"c30c30",
   12979 => x"c30c30",
   12980 => x"c30c30",
   12981 => x"c30c30",
   12982 => x"c30c28",
   12983 => x"b3cf3c",
   12984 => x"f3cf3c",
   12985 => x"f3cf3c",
   12986 => x"f3cf3c",
   12987 => x"f3cf3c",
   12988 => x"f3cf3c",
   12989 => x"f3cf3c",
   12990 => x"f3cf3c",
   12991 => x"f3cf3c",
   12992 => x"f3cf3c",
   12993 => x"f3cf3c",
   12994 => x"f3cf3c",
   12995 => x"f3cf3c",
   12996 => x"f3cf3c",
   12997 => x"f3cf3c",
   12998 => x"f3cf3c",
   12999 => x"f3cf3c",
   13000 => x"f3cf3c",
   13001 => x"f3cf3c",
   13002 => x"f3cf3c",
   13003 => x"f3cf3c",
   13004 => x"f3cf3c",
   13005 => x"f3cb0c",
   13006 => x"30c30c",
   13007 => x"30c30c",
   13008 => x"30c30c",
   13009 => x"30c30c",
   13010 => x"30c30c",
   13011 => x"30c30c",
   13012 => x"30c30c",
   13013 => x"30c30c",
   13014 => x"30c30c",
   13015 => x"30c30c",
   13016 => x"30c30c",
   13017 => x"30c30c",
   13018 => x"30c30c",
   13019 => x"30c30c",
   13020 => x"30c30c",
   13021 => x"30c30c",
   13022 => x"30c30c",
   13023 => x"30c30c",
   13024 => x"30c30c",
   13025 => x"30c30c",
   13026 => x"30c30c",
   13027 => x"30cbbf",
   13028 => x"ffffff",
   13029 => x"ffffff",
   13030 => x"ffffff",
   13031 => x"ffffff",
   13032 => x"ffffff",
   13033 => x"ffffff",
   13034 => x"ffffff",
   13035 => x"ffffff",
   13036 => x"ffffff",
   13037 => x"ffffff",
   13038 => x"ffffff",
   13039 => x"ffffff",
   13040 => x"ffffff",
   13041 => x"ffffff",
   13042 => x"ffffff",
   13043 => x"ffffff",
   13044 => x"ffffff",
   13045 => x"ffffff",
   13046 => x"ffffff",
   13047 => x"ffffff",
   13048 => x"ffffff",
   13049 => x"ffffff",
   13050 => x"ffffff",
   13051 => x"fea56a",
   13052 => x"ffffff",
   13053 => x"ffffff",
   13054 => x"ffffff",
   13055 => x"ffffff",
   13056 => x"ffffff",
   13057 => x"ffffff",
   13058 => x"ffffff",
   13059 => x"ffffff",
   13060 => x"ffffff",
   13061 => x"ffffff",
   13062 => x"ffffff",
   13063 => x"ffffff",
   13064 => x"ffffff",
   13065 => x"ffffff",
   13066 => x"ffffff",
   13067 => x"ffffff",
   13068 => x"ffffff",
   13069 => x"ffffff",
   13070 => x"ffffff",
   13071 => x"ffffff",
   13072 => x"ffffff",
   13073 => x"ffffff",
   13074 => x"ffffff",
   13075 => x"ffffff",
   13076 => x"ffffff",
   13077 => x"ffffff",
   13078 => x"ffffff",
   13079 => x"ffffff",
   13080 => x"ffffff",
   13081 => x"ffffff",
   13082 => x"ffffff",
   13083 => x"ffffff",
   13084 => x"ffffff",
   13085 => x"ffffff",
   13086 => x"ffffff",
   13087 => x"ffffff",
   13088 => x"ffffff",
   13089 => x"ffffff",
   13090 => x"ffffff",
   13091 => x"ffffff",
   13092 => x"ffffff",
   13093 => x"ffffff",
   13094 => x"ffffff",
   13095 => x"ffffff",
   13096 => x"ffffff",
   13097 => x"ffffff",
   13098 => x"ffffff",
   13099 => x"ffffff",
   13100 => x"ffffff",
   13101 => x"ffffff",
   13102 => x"ffffff",
   13103 => x"ffffff",
   13104 => x"ffffff",
   13105 => x"ffffff",
   13106 => x"ffffff",
   13107 => x"ffffff",
   13108 => x"ffffff",
   13109 => x"ffffff",
   13110 => x"ffffff",
   13111 => x"ffffff",
   13112 => x"ffffff",
   13113 => x"ffffff",
   13114 => x"ffffff",
   13115 => x"ffffff",
   13116 => x"ffffff",
   13117 => x"ffffff",
   13118 => x"ffffff",
   13119 => x"ffffff",
   13120 => x"ffffff",
   13121 => x"c30c30",
   13122 => x"c30c30",
   13123 => x"c30c30",
   13124 => x"c30c30",
   13125 => x"c30c30",
   13126 => x"c30c30",
   13127 => x"c30c30",
   13128 => x"c30c30",
   13129 => x"c30c30",
   13130 => x"c30c30",
   13131 => x"c30c30",
   13132 => x"c30c30",
   13133 => x"c30c30",
   13134 => x"c30c30",
   13135 => x"c30c30",
   13136 => x"c30c30",
   13137 => x"c30c30",
   13138 => x"c30c30",
   13139 => x"c30c30",
   13140 => x"c30c30",
   13141 => x"c30c30",
   13142 => x"c30c28",
   13143 => x"f3cf3c",
   13144 => x"f3cf3c",
   13145 => x"f3cf3c",
   13146 => x"f3cf3c",
   13147 => x"f3cf3c",
   13148 => x"f3cf3c",
   13149 => x"f3cf3c",
   13150 => x"f3cf3c",
   13151 => x"f3cf3c",
   13152 => x"f3cf3c",
   13153 => x"f3cf3c",
   13154 => x"f3cf3c",
   13155 => x"f3cf3c",
   13156 => x"f3cf3c",
   13157 => x"f3cf3c",
   13158 => x"f3cf3c",
   13159 => x"f3cf3c",
   13160 => x"f3cf3c",
   13161 => x"f3cf3c",
   13162 => x"f3cf3c",
   13163 => x"f3cf3c",
   13164 => x"f3cf3c",
   13165 => x"f3cb0c",
   13166 => x"30c30c",
   13167 => x"30c30c",
   13168 => x"30c30c",
   13169 => x"30c30c",
   13170 => x"30c30c",
   13171 => x"30c30c",
   13172 => x"30c30c",
   13173 => x"30c30c",
   13174 => x"30c30c",
   13175 => x"30c30c",
   13176 => x"30c30c",
   13177 => x"30c30c",
   13178 => x"30c30c",
   13179 => x"30c30c",
   13180 => x"30c30c",
   13181 => x"30c30c",
   13182 => x"30c30c",
   13183 => x"30c30c",
   13184 => x"30c30c",
   13185 => x"30c30c",
   13186 => x"30c30c",
   13187 => x"30c77f",
   13188 => x"ffffff",
   13189 => x"ffffff",
   13190 => x"ffffff",
   13191 => x"ffffff",
   13192 => x"ffffff",
   13193 => x"ffffff",
   13194 => x"ffffff",
   13195 => x"ffffff",
   13196 => x"ffffff",
   13197 => x"ffffff",
   13198 => x"ffffff",
   13199 => x"ffffff",
   13200 => x"ffffff",
   13201 => x"ffffff",
   13202 => x"ffffff",
   13203 => x"ffffff",
   13204 => x"ffffff",
   13205 => x"ffffff",
   13206 => x"ffffff",
   13207 => x"ffffff",
   13208 => x"ffffff",
   13209 => x"ffffff",
   13210 => x"ffffff",
   13211 => x"a95abf",
   13212 => x"ffffff",
   13213 => x"ffffff",
   13214 => x"ffffff",
   13215 => x"ffffff",
   13216 => x"ffffff",
   13217 => x"ffffff",
   13218 => x"ffffff",
   13219 => x"ffffff",
   13220 => x"ffffff",
   13221 => x"ffffff",
   13222 => x"ffffff",
   13223 => x"ffffff",
   13224 => x"ffffff",
   13225 => x"ffffff",
   13226 => x"ffffff",
   13227 => x"ffffff",
   13228 => x"ffffff",
   13229 => x"ffffff",
   13230 => x"ffffff",
   13231 => x"ffffff",
   13232 => x"ffffff",
   13233 => x"ffffff",
   13234 => x"ffffff",
   13235 => x"ffffff",
   13236 => x"ffffff",
   13237 => x"ffffff",
   13238 => x"ffffff",
   13239 => x"ffffff",
   13240 => x"ffffff",
   13241 => x"ffffff",
   13242 => x"ffffff",
   13243 => x"ffffff",
   13244 => x"ffffff",
   13245 => x"ffffff",
   13246 => x"ffffff",
   13247 => x"ffffff",
   13248 => x"ffffff",
   13249 => x"ffffff",
   13250 => x"ffffff",
   13251 => x"ffffff",
   13252 => x"ffffff",
   13253 => x"ffffff",
   13254 => x"ffffff",
   13255 => x"ffffff",
   13256 => x"ffffff",
   13257 => x"ffffff",
   13258 => x"ffffff",
   13259 => x"ffffff",
   13260 => x"ffffff",
   13261 => x"ffffff",
   13262 => x"ffffff",
   13263 => x"ffffff",
   13264 => x"ffffff",
   13265 => x"ffffff",
   13266 => x"ffffff",
   13267 => x"ffffff",
   13268 => x"ffffff",
   13269 => x"ffffff",
   13270 => x"ffffff",
   13271 => x"ffffff",
   13272 => x"ffffff",
   13273 => x"ffffff",
   13274 => x"ffffff",
   13275 => x"ffffff",
   13276 => x"ffffff",
   13277 => x"ffffff",
   13278 => x"ffffff",
   13279 => x"ffffff",
   13280 => x"fffffa",
   13281 => x"c30c30",
   13282 => x"c30c30",
   13283 => x"c30c30",
   13284 => x"c30c30",
   13285 => x"c30c30",
   13286 => x"c30c30",
   13287 => x"c30c30",
   13288 => x"c30c30",
   13289 => x"c30c30",
   13290 => x"c30c30",
   13291 => x"c30c30",
   13292 => x"c30c30",
   13293 => x"c30c30",
   13294 => x"c30c30",
   13295 => x"c30c30",
   13296 => x"c30c30",
   13297 => x"c30c30",
   13298 => x"c30c30",
   13299 => x"c30c30",
   13300 => x"c30c30",
   13301 => x"c30c30",
   13302 => x"c30928",
   13303 => x"f3cf3c",
   13304 => x"f3cf3c",
   13305 => x"f3cf3c",
   13306 => x"f3cf3c",
   13307 => x"f3cf3c",
   13308 => x"f3cf3c",
   13309 => x"f3cf3c",
   13310 => x"f3cf3c",
   13311 => x"f3cf3c",
   13312 => x"f3cf3c",
   13313 => x"f3cf3c",
   13314 => x"f3cf3c",
   13315 => x"f3cf3c",
   13316 => x"f3cf3c",
   13317 => x"f3cf3c",
   13318 => x"f3cf3c",
   13319 => x"f3cf3c",
   13320 => x"f3cf3c",
   13321 => x"f3cf3c",
   13322 => x"f3cf3c",
   13323 => x"f3cf3c",
   13324 => x"f3cf3c",
   13325 => x"f3cf1c",
   13326 => x"30c30c",
   13327 => x"30c30c",
   13328 => x"30c30c",
   13329 => x"30c30c",
   13330 => x"30c30c",
   13331 => x"30c30c",
   13332 => x"30c30c",
   13333 => x"30c30c",
   13334 => x"30c30c",
   13335 => x"30c30c",
   13336 => x"30c30c",
   13337 => x"30c30c",
   13338 => x"30c30c",
   13339 => x"30c30c",
   13340 => x"30c30c",
   13341 => x"30c30c",
   13342 => x"30c30c",
   13343 => x"30c30c",
   13344 => x"30c30c",
   13345 => x"30c30c",
   13346 => x"30c30c",
   13347 => x"30c77f",
   13348 => x"ffffff",
   13349 => x"ffffff",
   13350 => x"ffffff",
   13351 => x"ffffff",
   13352 => x"ffffff",
   13353 => x"ffffff",
   13354 => x"ffffff",
   13355 => x"ffffff",
   13356 => x"ffffff",
   13357 => x"ffffff",
   13358 => x"ffffff",
   13359 => x"ffffff",
   13360 => x"ffffff",
   13361 => x"ffffff",
   13362 => x"ffffff",
   13363 => x"ffffff",
   13364 => x"ffffff",
   13365 => x"ffffff",
   13366 => x"ffffff",
   13367 => x"ffffff",
   13368 => x"ffffff",
   13369 => x"ffffff",
   13370 => x"ffffea",
   13371 => x"56afff",
   13372 => x"ffffff",
   13373 => x"ffffff",
   13374 => x"ffffff",
   13375 => x"ffffff",
   13376 => x"ffffff",
   13377 => x"ffffff",
   13378 => x"ffffff",
   13379 => x"ffffff",
   13380 => x"ffffff",
   13381 => x"ffffff",
   13382 => x"ffffff",
   13383 => x"ffffff",
   13384 => x"ffffff",
   13385 => x"ffffff",
   13386 => x"ffffff",
   13387 => x"ffffff",
   13388 => x"ffffff",
   13389 => x"ffffff",
   13390 => x"ffffff",
   13391 => x"ffffff",
   13392 => x"ffffff",
   13393 => x"ffffff",
   13394 => x"ffffff",
   13395 => x"ffffff",
   13396 => x"ffffff",
   13397 => x"ffffff",
   13398 => x"ffffff",
   13399 => x"ffffff",
   13400 => x"ffffff",
   13401 => x"ffffff",
   13402 => x"ffffff",
   13403 => x"ffffff",
   13404 => x"ffffff",
   13405 => x"ffffff",
   13406 => x"ffffff",
   13407 => x"ffffff",
   13408 => x"ffffff",
   13409 => x"ffffff",
   13410 => x"ffffff",
   13411 => x"ffffff",
   13412 => x"ffffff",
   13413 => x"ffffff",
   13414 => x"ffffff",
   13415 => x"ffffff",
   13416 => x"ffffff",
   13417 => x"ffffff",
   13418 => x"ffffff",
   13419 => x"ffffff",
   13420 => x"ffffff",
   13421 => x"ffffff",
   13422 => x"ffffff",
   13423 => x"ffffff",
   13424 => x"ffffff",
   13425 => x"ffffff",
   13426 => x"ffffff",
   13427 => x"ffffff",
   13428 => x"ffffff",
   13429 => x"ffffff",
   13430 => x"ffffff",
   13431 => x"ffffff",
   13432 => x"ffffff",
   13433 => x"ffffff",
   13434 => x"ffffff",
   13435 => x"ffffff",
   13436 => x"ffffff",
   13437 => x"ffffff",
   13438 => x"ffffff",
   13439 => x"ffffff",
   13440 => x"fffff5",
   13441 => x"c30c30",
   13442 => x"c30c30",
   13443 => x"c30c30",
   13444 => x"c30c30",
   13445 => x"c30c30",
   13446 => x"c30c30",
   13447 => x"c30c30",
   13448 => x"c30c30",
   13449 => x"c30c30",
   13450 => x"c30c30",
   13451 => x"c30c30",
   13452 => x"c30c30",
   13453 => x"c30c30",
   13454 => x"c30c30",
   13455 => x"c30c30",
   13456 => x"c30c30",
   13457 => x"c30c30",
   13458 => x"c30c30",
   13459 => x"c30c30",
   13460 => x"c30c30",
   13461 => x"c30c30",
   13462 => x"c3092c",
   13463 => x"f3cf3c",
   13464 => x"f3cf3c",
   13465 => x"f3cf3c",
   13466 => x"f3cf3c",
   13467 => x"f3cf3c",
   13468 => x"f3cf3c",
   13469 => x"f3cf3c",
   13470 => x"f3cf3c",
   13471 => x"f3cf3c",
   13472 => x"f3cf3c",
   13473 => x"f3cf3c",
   13474 => x"f3cf3c",
   13475 => x"f3cf3c",
   13476 => x"f3cf3c",
   13477 => x"f3cf3c",
   13478 => x"f3cf3c",
   13479 => x"f3cf3c",
   13480 => x"f3cf3c",
   13481 => x"f3cf3c",
   13482 => x"f3cf3c",
   13483 => x"f3cf3c",
   13484 => x"f3cf3c",
   13485 => x"f3cf1c",
   13486 => x"30c30c",
   13487 => x"30c30c",
   13488 => x"30c30c",
   13489 => x"30c30c",
   13490 => x"30c30c",
   13491 => x"30c30c",
   13492 => x"30c30c",
   13493 => x"30c30c",
   13494 => x"30c30c",
   13495 => x"30c30c",
   13496 => x"30c30c",
   13497 => x"30c30c",
   13498 => x"30c30c",
   13499 => x"30c30c",
   13500 => x"30c30c",
   13501 => x"30c30c",
   13502 => x"30c30c",
   13503 => x"30c30c",
   13504 => x"30c30c",
   13505 => x"30c30c",
   13506 => x"30c30c",
   13507 => x"30c32e",
   13508 => x"ffffff",
   13509 => x"ffffff",
   13510 => x"ffffff",
   13511 => x"ffffff",
   13512 => x"ffffff",
   13513 => x"ffffff",
   13514 => x"ffffff",
   13515 => x"ffffff",
   13516 => x"ffffff",
   13517 => x"ffffff",
   13518 => x"ffffff",
   13519 => x"ffffff",
   13520 => x"ffffff",
   13521 => x"ffffff",
   13522 => x"ffffff",
   13523 => x"ffffff",
   13524 => x"ffffff",
   13525 => x"ffffff",
   13526 => x"ffffff",
   13527 => x"ffffff",
   13528 => x"ffffff",
   13529 => x"ffffff",
   13530 => x"fffa95",
   13531 => x"abffff",
   13532 => x"ffffff",
   13533 => x"ffffff",
   13534 => x"ffffff",
   13535 => x"ffffff",
   13536 => x"ffffff",
   13537 => x"ffffff",
   13538 => x"ffffff",
   13539 => x"ffffff",
   13540 => x"ffffff",
   13541 => x"ffffff",
   13542 => x"ffffff",
   13543 => x"ffffff",
   13544 => x"ffffff",
   13545 => x"ffffff",
   13546 => x"ffffff",
   13547 => x"ffffff",
   13548 => x"ffffff",
   13549 => x"ffffff",
   13550 => x"ffffff",
   13551 => x"ffffff",
   13552 => x"ffffff",
   13553 => x"ffffff",
   13554 => x"ffffff",
   13555 => x"ffffff",
   13556 => x"ffffff",
   13557 => x"ffffff",
   13558 => x"ffffff",
   13559 => x"ffffff",
   13560 => x"ffffff",
   13561 => x"ffffff",
   13562 => x"ffffff",
   13563 => x"ffffff",
   13564 => x"ffffff",
   13565 => x"ffffff",
   13566 => x"ffffff",
   13567 => x"ffffff",
   13568 => x"ffffff",
   13569 => x"ffffff",
   13570 => x"ffffff",
   13571 => x"ffffff",
   13572 => x"ffffff",
   13573 => x"ffffff",
   13574 => x"ffffff",
   13575 => x"ffffff",
   13576 => x"ffffff",
   13577 => x"ffffff",
   13578 => x"ffffff",
   13579 => x"ffffff",
   13580 => x"ffffff",
   13581 => x"ffffff",
   13582 => x"ffffff",
   13583 => x"ffffff",
   13584 => x"ffffff",
   13585 => x"ffffff",
   13586 => x"ffffff",
   13587 => x"ffffff",
   13588 => x"ffffff",
   13589 => x"ffffff",
   13590 => x"ffffff",
   13591 => x"ffffff",
   13592 => x"ffffff",
   13593 => x"ffffff",
   13594 => x"ffffff",
   13595 => x"ffffff",
   13596 => x"ffffff",
   13597 => x"ffffff",
   13598 => x"ffffff",
   13599 => x"ffffff",
   13600 => x"fffff5",
   13601 => x"c30c30",
   13602 => x"c30c30",
   13603 => x"c30c30",
   13604 => x"c30c30",
   13605 => x"c30c30",
   13606 => x"c30c30",
   13607 => x"c30c30",
   13608 => x"c30c30",
   13609 => x"c30c30",
   13610 => x"c30c30",
   13611 => x"c30c30",
   13612 => x"c30c30",
   13613 => x"c30c30",
   13614 => x"c30c30",
   13615 => x"c30c30",
   13616 => x"c30c30",
   13617 => x"c30c30",
   13618 => x"c30c30",
   13619 => x"c30c30",
   13620 => x"c30c30",
   13621 => x"c30c30",
   13622 => x"c30a2c",
   13623 => x"f3cf3c",
   13624 => x"f3cf3c",
   13625 => x"f3cf3c",
   13626 => x"f3cf3c",
   13627 => x"f3cf3c",
   13628 => x"f3cf3c",
   13629 => x"f3cf3c",
   13630 => x"f3cf3c",
   13631 => x"f3cf3c",
   13632 => x"f3cf3c",
   13633 => x"f3cf3c",
   13634 => x"f3cf3c",
   13635 => x"f3cf3c",
   13636 => x"f3cf3c",
   13637 => x"f3cf3c",
   13638 => x"f3cf3c",
   13639 => x"f3cf3c",
   13640 => x"f3cf3c",
   13641 => x"f3cf3c",
   13642 => x"f3cf3c",
   13643 => x"f3cf3c",
   13644 => x"f3cf3c",
   13645 => x"f3cf2c",
   13646 => x"30c30c",
   13647 => x"30c30c",
   13648 => x"30c30c",
   13649 => x"30c30c",
   13650 => x"30c30c",
   13651 => x"30c30c",
   13652 => x"30c30c",
   13653 => x"30c30c",
   13654 => x"30c30c",
   13655 => x"30c30c",
   13656 => x"30c30c",
   13657 => x"30c30c",
   13658 => x"30c30c",
   13659 => x"30c30c",
   13660 => x"30c30c",
   13661 => x"30c30c",
   13662 => x"30c30c",
   13663 => x"30c30c",
   13664 => x"30c30c",
   13665 => x"30c30c",
   13666 => x"30c30c",
   13667 => x"30c32e",
   13668 => x"ffffff",
   13669 => x"ffffff",
   13670 => x"ffffff",
   13671 => x"ffffff",
   13672 => x"ffffff",
   13673 => x"ffffff",
   13674 => x"ffffff",
   13675 => x"ffffff",
   13676 => x"ffffff",
   13677 => x"ffffff",
   13678 => x"ffffff",
   13679 => x"ffffff",
   13680 => x"ffffff",
   13681 => x"ffffff",
   13682 => x"ffffff",
   13683 => x"ffffff",
   13684 => x"ffffff",
   13685 => x"ffffff",
   13686 => x"ffffff",
   13687 => x"ffffff",
   13688 => x"ffffff",
   13689 => x"ffffff",
   13690 => x"fea56a",
   13691 => x"ffffff",
   13692 => x"ffffff",
   13693 => x"ffffff",
   13694 => x"ffffff",
   13695 => x"ffffff",
   13696 => x"ffffff",
   13697 => x"ffffff",
   13698 => x"ffffff",
   13699 => x"ffffff",
   13700 => x"ffffff",
   13701 => x"ffffff",
   13702 => x"ffffff",
   13703 => x"ffffff",
   13704 => x"ffffff",
   13705 => x"ffffff",
   13706 => x"ffffff",
   13707 => x"ffffff",
   13708 => x"ffffff",
   13709 => x"ffffff",
   13710 => x"ffffff",
   13711 => x"ffffff",
   13712 => x"ffffff",
   13713 => x"ffffff",
   13714 => x"ffffff",
   13715 => x"ffffff",
   13716 => x"ffffff",
   13717 => x"ffffff",
   13718 => x"ffffff",
   13719 => x"ffffff",
   13720 => x"ffffff",
   13721 => x"ffffff",
   13722 => x"ffffff",
   13723 => x"ffffff",
   13724 => x"ffffff",
   13725 => x"ffffff",
   13726 => x"ffffff",
   13727 => x"ffffff",
   13728 => x"ffffff",
   13729 => x"ffffff",
   13730 => x"ffffff",
   13731 => x"ffffff",
   13732 => x"ffffff",
   13733 => x"ffffff",
   13734 => x"ffffff",
   13735 => x"ffffff",
   13736 => x"ffffff",
   13737 => x"ffffff",
   13738 => x"ffffff",
   13739 => x"ffffff",
   13740 => x"ffffff",
   13741 => x"ffffff",
   13742 => x"ffffff",
   13743 => x"ffffff",
   13744 => x"ffffff",
   13745 => x"ffffff",
   13746 => x"ffffff",
   13747 => x"ffffff",
   13748 => x"ffffff",
   13749 => x"ffffff",
   13750 => x"ffffff",
   13751 => x"ffffff",
   13752 => x"ffffff",
   13753 => x"ffffff",
   13754 => x"ffffff",
   13755 => x"ffffff",
   13756 => x"ffffff",
   13757 => x"ffffff",
   13758 => x"ffffff",
   13759 => x"ffffff",
   13760 => x"fffff0",
   13761 => x"c30c30",
   13762 => x"c30c30",
   13763 => x"c30c30",
   13764 => x"c30c30",
   13765 => x"c30c30",
   13766 => x"c30c30",
   13767 => x"c30c30",
   13768 => x"c30c30",
   13769 => x"c30c30",
   13770 => x"c30c30",
   13771 => x"c30c30",
   13772 => x"c30c30",
   13773 => x"c30c30",
   13774 => x"c30c30",
   13775 => x"c30c30",
   13776 => x"c30c30",
   13777 => x"c30c30",
   13778 => x"c30c30",
   13779 => x"c30c30",
   13780 => x"c30c30",
   13781 => x"c30c30",
   13782 => x"c30a2c",
   13783 => x"f3cf3c",
   13784 => x"f3cf3c",
   13785 => x"f3cf3c",
   13786 => x"f3cf3c",
   13787 => x"f3cf3c",
   13788 => x"f3cf3c",
   13789 => x"f3cf3c",
   13790 => x"f3cf3c",
   13791 => x"f3cf3c",
   13792 => x"f3cf3c",
   13793 => x"f3cf3c",
   13794 => x"f3cf3c",
   13795 => x"f3cf3c",
   13796 => x"f3cf3c",
   13797 => x"f3cf3c",
   13798 => x"f3cf3c",
   13799 => x"f3cf3c",
   13800 => x"f3cf3c",
   13801 => x"f3cf3c",
   13802 => x"f3cf3c",
   13803 => x"f3cf3c",
   13804 => x"f3cf3c",
   13805 => x"f3cf2c",
   13806 => x"30c30c",
   13807 => x"30c30c",
   13808 => x"30c30c",
   13809 => x"30c30c",
   13810 => x"30c30c",
   13811 => x"30c30c",
   13812 => x"30c30c",
   13813 => x"30c30c",
   13814 => x"30c30c",
   13815 => x"30c30c",
   13816 => x"30c30c",
   13817 => x"30c30c",
   13818 => x"30c30c",
   13819 => x"30c30c",
   13820 => x"30c30c",
   13821 => x"30c30c",
   13822 => x"30c30c",
   13823 => x"30c30c",
   13824 => x"30c30c",
   13825 => x"30c30c",
   13826 => x"30c30c",
   13827 => x"30c32e",
   13828 => x"ffffff",
   13829 => x"ffffff",
   13830 => x"ffffff",
   13831 => x"ffffff",
   13832 => x"ffffff",
   13833 => x"ffffff",
   13834 => x"ffffff",
   13835 => x"ffffff",
   13836 => x"ffffff",
   13837 => x"ffffff",
   13838 => x"ffffff",
   13839 => x"ffffff",
   13840 => x"ffffff",
   13841 => x"ffffff",
   13842 => x"ffffff",
   13843 => x"ffffff",
   13844 => x"ffffff",
   13845 => x"ffffff",
   13846 => x"ffffff",
   13847 => x"ffffff",
   13848 => x"ffffff",
   13849 => x"ffffff",
   13850 => x"a95abf",
   13851 => x"ffffff",
   13852 => x"ffffff",
   13853 => x"ffffff",
   13854 => x"ffffff",
   13855 => x"ffffff",
   13856 => x"ffffff",
   13857 => x"ffffff",
   13858 => x"ffffff",
   13859 => x"ffffff",
   13860 => x"ffffff",
   13861 => x"ffffff",
   13862 => x"ffffff",
   13863 => x"ffffff",
   13864 => x"ffffff",
   13865 => x"ffffff",
   13866 => x"ffffff",
   13867 => x"ffffff",
   13868 => x"ffffff",
   13869 => x"ffffff",
   13870 => x"ffffff",
   13871 => x"ffffff",
   13872 => x"ffffff",
   13873 => x"ffffff",
   13874 => x"ffffff",
   13875 => x"ffffff",
   13876 => x"ffffff",
   13877 => x"ffffff",
   13878 => x"ffffff",
   13879 => x"ffffff",
   13880 => x"ffffff",
   13881 => x"ffffff",
   13882 => x"ffffff",
   13883 => x"ffffff",
   13884 => x"ffffff",
   13885 => x"ffffff",
   13886 => x"ffffff",
   13887 => x"ffffff",
   13888 => x"ffffff",
   13889 => x"ffffff",
   13890 => x"ffffff",
   13891 => x"ffffff",
   13892 => x"ffffff",
   13893 => x"ffffff",
   13894 => x"ffffff",
   13895 => x"ffffff",
   13896 => x"ffffff",
   13897 => x"ffffff",
   13898 => x"ffffff",
   13899 => x"ffffff",
   13900 => x"ffffff",
   13901 => x"ffffff",
   13902 => x"ffffff",
   13903 => x"ffffff",
   13904 => x"ffffff",
   13905 => x"ffffff",
   13906 => x"ffffff",
   13907 => x"ffffff",
   13908 => x"ffffff",
   13909 => x"ffffff",
   13910 => x"ffffff",
   13911 => x"ffffff",
   13912 => x"ffffff",
   13913 => x"ffffff",
   13914 => x"ffffff",
   13915 => x"ffffff",
   13916 => x"ffffff",
   13917 => x"ffffff",
   13918 => x"ffffff",
   13919 => x"ffffff",
   13920 => x"fffeb0",
   13921 => x"c30c30",
   13922 => x"c30c30",
   13923 => x"c30c30",
   13924 => x"c30c30",
   13925 => x"c30c30",
   13926 => x"c30c30",
   13927 => x"c30c30",
   13928 => x"c30c30",
   13929 => x"c30c30",
   13930 => x"c30c30",
   13931 => x"c30c30",
   13932 => x"c30c30",
   13933 => x"c30c30",
   13934 => x"c30c30",
   13935 => x"c30c30",
   13936 => x"c30c30",
   13937 => x"c30c30",
   13938 => x"c30c30",
   13939 => x"c30c30",
   13940 => x"c30c30",
   13941 => x"c30c30",
   13942 => x"c30a3c",
   13943 => x"f3cf3c",
   13944 => x"f3cf3c",
   13945 => x"f3cf3c",
   13946 => x"f3cf3c",
   13947 => x"f3cf3c",
   13948 => x"f3cf3c",
   13949 => x"f3cf3c",
   13950 => x"f3cf3c",
   13951 => x"f3cf3c",
   13952 => x"f3cf3c",
   13953 => x"f3cf3c",
   13954 => x"f3cf3c",
   13955 => x"f3cf3c",
   13956 => x"f3cf3c",
   13957 => x"f3cf3c",
   13958 => x"f3cf3c",
   13959 => x"f3cf3c",
   13960 => x"f3cf3c",
   13961 => x"f3cf3c",
   13962 => x"f3cf3c",
   13963 => x"f3cf3c",
   13964 => x"f3cf3c",
   13965 => x"f3cf3c",
   13966 => x"30c30c",
   13967 => x"30c30c",
   13968 => x"30c30c",
   13969 => x"30c30c",
   13970 => x"30c30c",
   13971 => x"30c30c",
   13972 => x"30c30c",
   13973 => x"30c30c",
   13974 => x"30c30c",
   13975 => x"30c30c",
   13976 => x"30c30c",
   13977 => x"30c30c",
   13978 => x"30c30c",
   13979 => x"30c30c",
   13980 => x"30c30c",
   13981 => x"30c30c",
   13982 => x"30c30c",
   13983 => x"30c30c",
   13984 => x"30c30c",
   13985 => x"30c30c",
   13986 => x"30c30c",
   13987 => x"30c31d",
   13988 => x"ffffff",
   13989 => x"ffffff",
   13990 => x"ffffff",
   13991 => x"ffffff",
   13992 => x"ffffff",
   13993 => x"ffffff",
   13994 => x"ffffff",
   13995 => x"ffffff",
   13996 => x"ffffff",
   13997 => x"ffffff",
   13998 => x"ffffff",
   13999 => x"ffffff",
   14000 => x"ffffff",
   14001 => x"ffffff",
   14002 => x"ffffff",
   14003 => x"ffffff",
   14004 => x"ffffff",
   14005 => x"ffffff",
   14006 => x"ffffff",
   14007 => x"ffffff",
   14008 => x"ffffff",
   14009 => x"ffffea",
   14010 => x"56afff",
   14011 => x"ffffff",
   14012 => x"ffffff",
   14013 => x"ffffff",
   14014 => x"ffffff",
   14015 => x"ffffff",
   14016 => x"ffffff",
   14017 => x"ffffff",
   14018 => x"ffffff",
   14019 => x"ffffff",
   14020 => x"ffffff",
   14021 => x"ffffff",
   14022 => x"ffffff",
   14023 => x"ffffff",
   14024 => x"ffffff",
   14025 => x"ffffff",
   14026 => x"ffffff",
   14027 => x"ffffff",
   14028 => x"ffffff",
   14029 => x"ffffff",
   14030 => x"ffffff",
   14031 => x"ffffff",
   14032 => x"ffffff",
   14033 => x"ffffff",
   14034 => x"ffffff",
   14035 => x"ffffff",
   14036 => x"ffffff",
   14037 => x"ffffff",
   14038 => x"ffffff",
   14039 => x"ffffff",
   14040 => x"ffffff",
   14041 => x"ffffff",
   14042 => x"ffffff",
   14043 => x"ffffff",
   14044 => x"ffffff",
   14045 => x"ffffff",
   14046 => x"ffffff",
   14047 => x"ffffff",
   14048 => x"ffffff",
   14049 => x"ffffff",
   14050 => x"ffffff",
   14051 => x"ffffff",
   14052 => x"ffffff",
   14053 => x"ffffff",
   14054 => x"ffffff",
   14055 => x"ffffff",
   14056 => x"ffffff",
   14057 => x"ffffff",
   14058 => x"ffffff",
   14059 => x"ffffff",
   14060 => x"ffffff",
   14061 => x"ffffff",
   14062 => x"ffffff",
   14063 => x"ffffff",
   14064 => x"ffffff",
   14065 => x"ffffff",
   14066 => x"ffffff",
   14067 => x"ffffff",
   14068 => x"ffffff",
   14069 => x"ffffff",
   14070 => x"ffffff",
   14071 => x"ffffff",
   14072 => x"ffffff",
   14073 => x"ffffff",
   14074 => x"ffffff",
   14075 => x"ffffff",
   14076 => x"ffffff",
   14077 => x"ffffff",
   14078 => x"ffffff",
   14079 => x"ffffff",
   14080 => x"fffeb0",
   14081 => x"c30c30",
   14082 => x"c30c30",
   14083 => x"c30c30",
   14084 => x"c30c30",
   14085 => x"c30c30",
   14086 => x"c30c30",
   14087 => x"c30c30",
   14088 => x"c30c30",
   14089 => x"c30c30",
   14090 => x"c30c30",
   14091 => x"c30c30",
   14092 => x"c30c30",
   14093 => x"c30c30",
   14094 => x"c30c30",
   14095 => x"c30c30",
   14096 => x"c30c30",
   14097 => x"c30c30",
   14098 => x"c30c30",
   14099 => x"c30c30",
   14100 => x"c30c30",
   14101 => x"c30c30",
   14102 => x"c24a3c",
   14103 => x"f3cf3c",
   14104 => x"f3cf3c",
   14105 => x"f3cf3c",
   14106 => x"f3cf3c",
   14107 => x"f3cf3c",
   14108 => x"f3cf3c",
   14109 => x"f3cf3c",
   14110 => x"f3cf3c",
   14111 => x"f3cf3c",
   14112 => x"f3cf3c",
   14113 => x"f3cf3c",
   14114 => x"f3cf3c",
   14115 => x"f3cf3c",
   14116 => x"f3cf3c",
   14117 => x"f3cf3c",
   14118 => x"f3cf3c",
   14119 => x"f3cf3c",
   14120 => x"f3cf3c",
   14121 => x"f3cf3c",
   14122 => x"f3cf3c",
   14123 => x"f3cf3c",
   14124 => x"f3cf3c",
   14125 => x"f3cf3c",
   14126 => x"70c30c",
   14127 => x"30c30c",
   14128 => x"30c30c",
   14129 => x"30c30c",
   14130 => x"30c30c",
   14131 => x"30c30c",
   14132 => x"30c30c",
   14133 => x"30c30c",
   14134 => x"30c30c",
   14135 => x"30c30c",
   14136 => x"30c30c",
   14137 => x"30c30c",
   14138 => x"30c30c",
   14139 => x"30c30c",
   14140 => x"30c30c",
   14141 => x"30c30c",
   14142 => x"30c30c",
   14143 => x"30c30c",
   14144 => x"30c30c",
   14145 => x"30c30c",
   14146 => x"30c30c",
   14147 => x"30c31d",
   14148 => x"ffffff",
   14149 => x"ffffff",
   14150 => x"ffffff",
   14151 => x"ffffff",
   14152 => x"ffffff",
   14153 => x"ffffff",
   14154 => x"ffffff",
   14155 => x"ffffff",
   14156 => x"ffffff",
   14157 => x"ffffff",
   14158 => x"ffffff",
   14159 => x"ffffff",
   14160 => x"ffffff",
   14161 => x"ffffff",
   14162 => x"ffffff",
   14163 => x"ffffff",
   14164 => x"ffffff",
   14165 => x"ffffff",
   14166 => x"ffffff",
   14167 => x"ffffff",
   14168 => x"ffffff",
   14169 => x"fffa95",
   14170 => x"abffff",
   14171 => x"ffffff",
   14172 => x"ffffff",
   14173 => x"ffffff",
   14174 => x"ffffff",
   14175 => x"ffffff",
   14176 => x"ffffff",
   14177 => x"ffffff",
   14178 => x"ffffff",
   14179 => x"ffffff",
   14180 => x"ffffff",
   14181 => x"ffffff",
   14182 => x"ffffff",
   14183 => x"ffffff",
   14184 => x"ffffff",
   14185 => x"ffffff",
   14186 => x"ffffff",
   14187 => x"ffffff",
   14188 => x"ffffff",
   14189 => x"ffffff",
   14190 => x"ffffff",
   14191 => x"ffffff",
   14192 => x"ffffff",
   14193 => x"ffffff",
   14194 => x"ffffff",
   14195 => x"ffffff",
   14196 => x"ffffff",
   14197 => x"ffffff",
   14198 => x"ffffff",
   14199 => x"ffffff",
   14200 => x"ffffff",
   14201 => x"ffffff",
   14202 => x"ffffff",
   14203 => x"ffffff",
   14204 => x"ffffff",
   14205 => x"ffffff",
   14206 => x"ffffff",
   14207 => x"ffffff",
   14208 => x"ffffff",
   14209 => x"ffffff",
   14210 => x"ffffff",
   14211 => x"ffffff",
   14212 => x"ffffff",
   14213 => x"ffffff",
   14214 => x"ffffff",
   14215 => x"ffffff",
   14216 => x"ffffff",
   14217 => x"ffffff",
   14218 => x"ffffff",
   14219 => x"ffffff",
   14220 => x"ffffff",
   14221 => x"ffffff",
   14222 => x"ffffff",
   14223 => x"ffffff",
   14224 => x"ffffff",
   14225 => x"ffffff",
   14226 => x"ffffff",
   14227 => x"ffffff",
   14228 => x"ffffff",
   14229 => x"ffffff",
   14230 => x"ffffff",
   14231 => x"ffffff",
   14232 => x"ffffff",
   14233 => x"ffffff",
   14234 => x"ffffff",
   14235 => x"ffffff",
   14236 => x"ffffff",
   14237 => x"ffffff",
   14238 => x"ffffff",
   14239 => x"ffffff",
   14240 => x"fffeb0",
   14241 => x"c30c30",
   14242 => x"c30c30",
   14243 => x"c30c30",
   14244 => x"c30c30",
   14245 => x"c30c30",
   14246 => x"c30c30",
   14247 => x"c30c30",
   14248 => x"c30c30",
   14249 => x"c30c30",
   14250 => x"c30c30",
   14251 => x"c30c30",
   14252 => x"c30c30",
   14253 => x"c30c30",
   14254 => x"c30c30",
   14255 => x"c30c30",
   14256 => x"c30c30",
   14257 => x"c30c30",
   14258 => x"c30c30",
   14259 => x"c30c30",
   14260 => x"c30c30",
   14261 => x"c30c30",
   14262 => x"c24b3c",
   14263 => x"f3cf3c",
   14264 => x"f3cf3c",
   14265 => x"f3cf3c",
   14266 => x"f3cf3c",
   14267 => x"f3cf3c",
   14268 => x"f3cf3c",
   14269 => x"f3cf3c",
   14270 => x"f3cf3c",
   14271 => x"f3cf3c",
   14272 => x"f3cf3c",
   14273 => x"f3cf3c",
   14274 => x"f3cf3c",
   14275 => x"f3cf3c",
   14276 => x"f3cf3c",
   14277 => x"f3cf3c",
   14278 => x"f3cf3c",
   14279 => x"f3cf3c",
   14280 => x"f3cf3c",
   14281 => x"f3cf3c",
   14282 => x"f3cf3c",
   14283 => x"f3cf3c",
   14284 => x"f3cf3c",
   14285 => x"f3cf3c",
   14286 => x"70c30c",
   14287 => x"30c30c",
   14288 => x"30c30c",
   14289 => x"30c30c",
   14290 => x"30c30c",
   14291 => x"30c30c",
   14292 => x"30c30c",
   14293 => x"30c30c",
   14294 => x"30c30c",
   14295 => x"30c30c",
   14296 => x"30c30c",
   14297 => x"30c30c",
   14298 => x"30c30c",
   14299 => x"30c30c",
   14300 => x"30c30c",
   14301 => x"30c30c",
   14302 => x"30c30c",
   14303 => x"30c30c",
   14304 => x"30c30c",
   14305 => x"30c30c",
   14306 => x"30c30c",
   14307 => x"30c30c",
   14308 => x"bbffff",
   14309 => x"ffffff",
   14310 => x"ffffff",
   14311 => x"ffffff",
   14312 => x"ffffff",
   14313 => x"ffffff",
   14314 => x"ffffff",
   14315 => x"ffffff",
   14316 => x"ffffff",
   14317 => x"ffffff",
   14318 => x"ffffff",
   14319 => x"ffffff",
   14320 => x"ffffff",
   14321 => x"ffffff",
   14322 => x"ffffff",
   14323 => x"ffffff",
   14324 => x"ffffff",
   14325 => x"ffffff",
   14326 => x"ffffff",
   14327 => x"ffffff",
   14328 => x"ffffff",
   14329 => x"fea56a",
   14330 => x"ffffff",
   14331 => x"ffffff",
   14332 => x"ffffff",
   14333 => x"ffffff",
   14334 => x"ffffff",
   14335 => x"ffffff",
   14336 => x"ffffff",
   14337 => x"ffffff",
   14338 => x"ffffff",
   14339 => x"ffffff",
   14340 => x"ffffff",
   14341 => x"ffffff",
   14342 => x"ffffff",
   14343 => x"ffffff",
   14344 => x"ffffff",
   14345 => x"ffffff",
   14346 => x"ffffff",
   14347 => x"ffffff",
   14348 => x"ffffff",
   14349 => x"ffffff",
   14350 => x"ffffff",
   14351 => x"ffffff",
   14352 => x"ffffff",
   14353 => x"ffffff",
   14354 => x"ffffff",
   14355 => x"ffffff",
   14356 => x"ffffff",
   14357 => x"ffffff",
   14358 => x"ffffff",
   14359 => x"ffffff",
   14360 => x"ffffff",
   14361 => x"ffffff",
   14362 => x"ffffff",
   14363 => x"ffffff",
   14364 => x"ffffff",
   14365 => x"ffffff",
   14366 => x"ffffff",
   14367 => x"ffffff",
   14368 => x"ffffff",
   14369 => x"ffffff",
   14370 => x"ffffff",
   14371 => x"ffffff",
   14372 => x"ffffff",
   14373 => x"ffffff",
   14374 => x"ffffff",
   14375 => x"ffffff",
   14376 => x"ffffff",
   14377 => x"ffffff",
   14378 => x"ffffff",
   14379 => x"ffffff",
   14380 => x"ffffff",
   14381 => x"ffffff",
   14382 => x"ffffff",
   14383 => x"ffffff",
   14384 => x"ffffff",
   14385 => x"ffffff",
   14386 => x"ffffff",
   14387 => x"ffffff",
   14388 => x"ffffff",
   14389 => x"ffffff",
   14390 => x"ffffff",
   14391 => x"ffffff",
   14392 => x"ffffff",
   14393 => x"ffffff",
   14394 => x"ffffff",
   14395 => x"ffffff",
   14396 => x"ffffff",
   14397 => x"ffffff",
   14398 => x"ffffff",
   14399 => x"ffffff",
   14400 => x"fffd70",
   14401 => x"c30c30",
   14402 => x"c30c30",
   14403 => x"c30c30",
   14404 => x"c30c30",
   14405 => x"c30c30",
   14406 => x"c30c30",
   14407 => x"c30c30",
   14408 => x"c30c30",
   14409 => x"c30c30",
   14410 => x"c30c30",
   14411 => x"c30c30",
   14412 => x"c30c30",
   14413 => x"c30c30",
   14414 => x"c30c30",
   14415 => x"c30c30",
   14416 => x"c30c30",
   14417 => x"c30c30",
   14418 => x"c30c30",
   14419 => x"c30c30",
   14420 => x"c30c30",
   14421 => x"c30c30",
   14422 => x"c24b3c",
   14423 => x"f3cf3c",
   14424 => x"f3cf3c",
   14425 => x"f3cf3c",
   14426 => x"f3cf3c",
   14427 => x"f3cf3c",
   14428 => x"f3cf3c",
   14429 => x"f3cf3c",
   14430 => x"f3cf3c",
   14431 => x"f3cf3c",
   14432 => x"f3cf3c",
   14433 => x"f3cf3c",
   14434 => x"f3cf3c",
   14435 => x"f3cf3c",
   14436 => x"f3cf3c",
   14437 => x"f3cf3c",
   14438 => x"f3cf3c",
   14439 => x"f3cf3c",
   14440 => x"f3cf3c",
   14441 => x"f3cf3c",
   14442 => x"f3cf3c",
   14443 => x"f3cf3c",
   14444 => x"f3cf3c",
   14445 => x"f3cf3c",
   14446 => x"70c30c",
   14447 => x"30c30c",
   14448 => x"30c30c",
   14449 => x"30c30c",
   14450 => x"30c30c",
   14451 => x"30c30c",
   14452 => x"30c30c",
   14453 => x"30c30c",
   14454 => x"30c30c",
   14455 => x"30c30c",
   14456 => x"30c30c",
   14457 => x"30c30c",
   14458 => x"30c30c",
   14459 => x"30c30c",
   14460 => x"30c30c",
   14461 => x"30c30c",
   14462 => x"30c30c",
   14463 => x"30c30c",
   14464 => x"30c30c",
   14465 => x"30c30c",
   14466 => x"30c30c",
   14467 => x"30c30c",
   14468 => x"bbffff",
   14469 => x"ffffff",
   14470 => x"ffffff",
   14471 => x"ffffff",
   14472 => x"ffffff",
   14473 => x"ffffff",
   14474 => x"ffffff",
   14475 => x"ffffff",
   14476 => x"ffffff",
   14477 => x"ffffff",
   14478 => x"ffffff",
   14479 => x"ffffff",
   14480 => x"ffffff",
   14481 => x"ffffff",
   14482 => x"ffffff",
   14483 => x"ffffff",
   14484 => x"ffffff",
   14485 => x"ffffff",
   14486 => x"ffffff",
   14487 => x"ffffff",
   14488 => x"ffffff",
   14489 => x"a95abf",
   14490 => x"ffffff",
   14491 => x"ffffff",
   14492 => x"ffffff",
   14493 => x"ffffff",
   14494 => x"ffffff",
   14495 => x"ffffff",
   14496 => x"ffffff",
   14497 => x"ffffff",
   14498 => x"ffffff",
   14499 => x"ffffff",
   14500 => x"ffffff",
   14501 => x"ffffff",
   14502 => x"ffffff",
   14503 => x"ffffff",
   14504 => x"ffffff",
   14505 => x"ffffff",
   14506 => x"ffffff",
   14507 => x"ffffff",
   14508 => x"ffffff",
   14509 => x"ffffff",
   14510 => x"ffffff",
   14511 => x"ffffff",
   14512 => x"ffffff",
   14513 => x"ffffff",
   14514 => x"ffffff",
   14515 => x"ffffff",
   14516 => x"ffffff",
   14517 => x"ffffff",
   14518 => x"ffffff",
   14519 => x"ffffff",
   14520 => x"ffffff",
   14521 => x"ffffff",
   14522 => x"ffffff",
   14523 => x"ffffff",
   14524 => x"ffffff",
   14525 => x"ffffff",
   14526 => x"ffffff",
   14527 => x"ffffff",
   14528 => x"ffffff",
   14529 => x"ffffff",
   14530 => x"ffffff",
   14531 => x"ffffff",
   14532 => x"ffffff",
   14533 => x"ffffff",
   14534 => x"ffffff",
   14535 => x"ffffff",
   14536 => x"ffffff",
   14537 => x"ffffff",
   14538 => x"ffffff",
   14539 => x"ffffff",
   14540 => x"ffffff",
   14541 => x"ffffff",
   14542 => x"ffffff",
   14543 => x"ffffff",
   14544 => x"ffffff",
   14545 => x"ffffff",
   14546 => x"ffffff",
   14547 => x"ffffff",
   14548 => x"ffffff",
   14549 => x"ffffff",
   14550 => x"ffffff",
   14551 => x"ffffff",
   14552 => x"ffffff",
   14553 => x"ffffff",
   14554 => x"ffffff",
   14555 => x"ffffff",
   14556 => x"ffffff",
   14557 => x"ffffff",
   14558 => x"ffffff",
   14559 => x"ffffff",
   14560 => x"fffd70",
   14561 => x"c30c30",
   14562 => x"c30c30",
   14563 => x"c30c30",
   14564 => x"c30c30",
   14565 => x"c30c30",
   14566 => x"c30c30",
   14567 => x"c30c30",
   14568 => x"c30c30",
   14569 => x"c30c30",
   14570 => x"c30c30",
   14571 => x"c30c30",
   14572 => x"c30c30",
   14573 => x"c30c30",
   14574 => x"c30c30",
   14575 => x"c30c30",
   14576 => x"c30c30",
   14577 => x"c30c30",
   14578 => x"c30c30",
   14579 => x"c30c30",
   14580 => x"c30c30",
   14581 => x"c30c30",
   14582 => x"c28b3c",
   14583 => x"f3cf3c",
   14584 => x"f3cf3c",
   14585 => x"f3cf3c",
   14586 => x"f3cf3c",
   14587 => x"f3cf3c",
   14588 => x"f3cf3c",
   14589 => x"f3cf3c",
   14590 => x"f3cf3c",
   14591 => x"f3cf3c",
   14592 => x"f3cf3c",
   14593 => x"f3cf3c",
   14594 => x"f3cf3c",
   14595 => x"f3cf3c",
   14596 => x"f3cf3c",
   14597 => x"f3cf3c",
   14598 => x"f3cf3c",
   14599 => x"f3cf3c",
   14600 => x"f3cf3c",
   14601 => x"f3cf3c",
   14602 => x"f3cf3c",
   14603 => x"f3cf3c",
   14604 => x"f3cf3c",
   14605 => x"f3cf3c",
   14606 => x"70c30c",
   14607 => x"30c30c",
   14608 => x"30c30c",
   14609 => x"30c30c",
   14610 => x"30c30c",
   14611 => x"30c30c",
   14612 => x"30c30c",
   14613 => x"30c30c",
   14614 => x"30c30c",
   14615 => x"30c30c",
   14616 => x"30c30c",
   14617 => x"30c30c",
   14618 => x"30c30c",
   14619 => x"30c30c",
   14620 => x"30c30c",
   14621 => x"30c30c",
   14622 => x"30c30c",
   14623 => x"30c30c",
   14624 => x"30c30c",
   14625 => x"30c30c",
   14626 => x"30c30c",
   14627 => x"30c30c",
   14628 => x"bbffff",
   14629 => x"ffffff",
   14630 => x"ffffff",
   14631 => x"ffffff",
   14632 => x"ffffff",
   14633 => x"ffffff",
   14634 => x"ffffff",
   14635 => x"ffffff",
   14636 => x"ffffff",
   14637 => x"ffffff",
   14638 => x"ffffff",
   14639 => x"ffffff",
   14640 => x"ffffff",
   14641 => x"ffffff",
   14642 => x"ffffff",
   14643 => x"ffffff",
   14644 => x"ffffff",
   14645 => x"ffffff",
   14646 => x"ffffff",
   14647 => x"ffffff",
   14648 => x"ffffea",
   14649 => x"56afff",
   14650 => x"ffffff",
   14651 => x"ffffff",
   14652 => x"ffffff",
   14653 => x"ffffff",
   14654 => x"ffffff",
   14655 => x"ffffff",
   14656 => x"ffffff",
   14657 => x"ffffff",
   14658 => x"ffffff",
   14659 => x"ffffff",
   14660 => x"ffffff",
   14661 => x"ffffff",
   14662 => x"ffffff",
   14663 => x"ffffff",
   14664 => x"ffffff",
   14665 => x"ffffff",
   14666 => x"ffffff",
   14667 => x"ffffff",
   14668 => x"ffffff",
   14669 => x"ffffff",
   14670 => x"ffffff",
   14671 => x"ffffff",
   14672 => x"ffffff",
   14673 => x"ffffff",
   14674 => x"ffffff",
   14675 => x"ffffff",
   14676 => x"ffffff",
   14677 => x"ffffff",
   14678 => x"ffffff",
   14679 => x"ffffff",
   14680 => x"ffffff",
   14681 => x"ffffff",
   14682 => x"ffffff",
   14683 => x"ffffff",
   14684 => x"ffffff",
   14685 => x"ffffff",
   14686 => x"ffffff",
   14687 => x"ffffff",
   14688 => x"ffffff",
   14689 => x"ffffff",
   14690 => x"ffffff",
   14691 => x"ffffff",
   14692 => x"ffffff",
   14693 => x"ffffff",
   14694 => x"ffffff",
   14695 => x"ffffff",
   14696 => x"ffffff",
   14697 => x"ffffff",
   14698 => x"ffffff",
   14699 => x"ffffff",
   14700 => x"ffffff",
   14701 => x"ffffff",
   14702 => x"ffffff",
   14703 => x"ffffff",
   14704 => x"ffffff",
   14705 => x"ffffff",
   14706 => x"ffffff",
   14707 => x"ffffff",
   14708 => x"ffffff",
   14709 => x"ffffff",
   14710 => x"ffffff",
   14711 => x"ffffff",
   14712 => x"ffffff",
   14713 => x"ffffff",
   14714 => x"ffffff",
   14715 => x"ffffff",
   14716 => x"ffffff",
   14717 => x"ffffff",
   14718 => x"ffffff",
   14719 => x"ffffff",
   14720 => x"fffd70",
   14721 => x"c30c30",
   14722 => x"c30c30",
   14723 => x"c30c30",
   14724 => x"c30c30",
   14725 => x"c30c30",
   14726 => x"c30c30",
   14727 => x"c30c30",
   14728 => x"c30c30",
   14729 => x"c30c30",
   14730 => x"c30c30",
   14731 => x"c30c30",
   14732 => x"c30c30",
   14733 => x"c30c30",
   14734 => x"c30c30",
   14735 => x"c30c30",
   14736 => x"c30c30",
   14737 => x"c30c30",
   14738 => x"c30c30",
   14739 => x"c30c30",
   14740 => x"c30c30",
   14741 => x"c30c30",
   14742 => x"c28b3c",
   14743 => x"f3cf3c",
   14744 => x"f3cf3c",
   14745 => x"f3cf3c",
   14746 => x"f3cf3c",
   14747 => x"f3cf3c",
   14748 => x"f3cf3c",
   14749 => x"f3cf3c",
   14750 => x"f3cf3c",
   14751 => x"f3cf3c",
   14752 => x"f3cf3c",
   14753 => x"f3cf3c",
   14754 => x"f3cf3c",
   14755 => x"f3cf3c",
   14756 => x"f3cf3c",
   14757 => x"f3cf3c",
   14758 => x"f3cf3c",
   14759 => x"f3cf3c",
   14760 => x"f3cf3c",
   14761 => x"f3cf3c",
   14762 => x"f3cf3c",
   14763 => x"f3cf3c",
   14764 => x"f3cf3c",
   14765 => x"f3cf3c",
   14766 => x"b0c30c",
   14767 => x"30c30c",
   14768 => x"30c30c",
   14769 => x"30c30c",
   14770 => x"30c30c",
   14771 => x"30c30c",
   14772 => x"30c30c",
   14773 => x"30c30c",
   14774 => x"30c30c",
   14775 => x"30c30c",
   14776 => x"30c30c",
   14777 => x"30c30c",
   14778 => x"30c30c",
   14779 => x"30c30c",
   14780 => x"30c30c",
   14781 => x"30c30c",
   14782 => x"30c30c",
   14783 => x"30c30c",
   14784 => x"30c30c",
   14785 => x"30c30c",
   14786 => x"30c30c",
   14787 => x"30c30c",
   14788 => x"bbffff",
   14789 => x"ffffff",
   14790 => x"ffffff",
   14791 => x"ffffff",
   14792 => x"ffffff",
   14793 => x"ffffff",
   14794 => x"ffffff",
   14795 => x"ffffff",
   14796 => x"ffffff",
   14797 => x"ffffff",
   14798 => x"ffffff",
   14799 => x"ffffff",
   14800 => x"ffffff",
   14801 => x"ffffff",
   14802 => x"ffffff",
   14803 => x"ffffff",
   14804 => x"ffffff",
   14805 => x"ffffff",
   14806 => x"ffffff",
   14807 => x"ffffff",
   14808 => x"fffa95",
   14809 => x"abffff",
   14810 => x"ffffff",
   14811 => x"ffffff",
   14812 => x"ffffff",
   14813 => x"ffffff",
   14814 => x"ffffff",
   14815 => x"ffffff",
   14816 => x"ffffff",
   14817 => x"ffffff",
   14818 => x"ffffff",
   14819 => x"ffffff",
   14820 => x"ffffff",
   14821 => x"ffffff",
   14822 => x"ffffff",
   14823 => x"ffffff",
   14824 => x"ffffff",
   14825 => x"ffffff",
   14826 => x"ffffff",
   14827 => x"ffffff",
   14828 => x"ffffff",
   14829 => x"ffffff",
   14830 => x"ffffff",
   14831 => x"ffffff",
   14832 => x"ffffff",
   14833 => x"ffffff",
   14834 => x"ffffff",
   14835 => x"ffffff",
   14836 => x"ffffff",
   14837 => x"ffffff",
   14838 => x"ffffff",
   14839 => x"ffffff",
   14840 => x"ffffff",
   14841 => x"ffffff",
   14842 => x"ffffff",
   14843 => x"ffffff",
   14844 => x"ffffff",
   14845 => x"ffffff",
   14846 => x"ffffff",
   14847 => x"ffffff",
   14848 => x"ffffff",
   14849 => x"ffffff",
   14850 => x"ffffff",
   14851 => x"ffffff",
   14852 => x"ffffff",
   14853 => x"ffffff",
   14854 => x"ffffff",
   14855 => x"ffffff",
   14856 => x"ffffff",
   14857 => x"ffffff",
   14858 => x"ffffff",
   14859 => x"ffffff",
   14860 => x"ffffff",
   14861 => x"ffffff",
   14862 => x"ffffff",
   14863 => x"ffffff",
   14864 => x"ffffff",
   14865 => x"ffffff",
   14866 => x"ffffff",
   14867 => x"ffffff",
   14868 => x"ffffff",
   14869 => x"ffffff",
   14870 => x"ffffff",
   14871 => x"ffffff",
   14872 => x"ffffff",
   14873 => x"ffffff",
   14874 => x"ffffff",
   14875 => x"ffffff",
   14876 => x"ffffff",
   14877 => x"ffffff",
   14878 => x"ffffff",
   14879 => x"ffffff",
   14880 => x"fffc30",
   14881 => x"c30c30",
   14882 => x"c30c30",
   14883 => x"c30c30",
   14884 => x"c30c30",
   14885 => x"c30c30",
   14886 => x"c30c30",
   14887 => x"c30c30",
   14888 => x"c30c30",
   14889 => x"c30c30",
   14890 => x"c30c30",
   14891 => x"c30c30",
   14892 => x"c30c30",
   14893 => x"c30c30",
   14894 => x"c30c30",
   14895 => x"c30c30",
   14896 => x"c30c30",
   14897 => x"c30c30",
   14898 => x"c30c30",
   14899 => x"c30c30",
   14900 => x"c30c30",
   14901 => x"c30c30",
   14902 => x"c28b3c",
   14903 => x"f3cf3c",
   14904 => x"f3cf3c",
   14905 => x"f3cf3c",
   14906 => x"f3cf3c",
   14907 => x"f3cf3c",
   14908 => x"f3cf3c",
   14909 => x"f3cf3c",
   14910 => x"f3cf3c",
   14911 => x"f3cf3c",
   14912 => x"f3cf3c",
   14913 => x"f3cf3c",
   14914 => x"f3cf3c",
   14915 => x"f3cf3c",
   14916 => x"f3cf3c",
   14917 => x"f3cf3c",
   14918 => x"f3cf3c",
   14919 => x"f3cf3c",
   14920 => x"f3cf3c",
   14921 => x"f3cf3c",
   14922 => x"f3cf3c",
   14923 => x"f3cf3c",
   14924 => x"f3cf3c",
   14925 => x"f3cf3c",
   14926 => x"b0c30c",
   14927 => x"30c30c",
   14928 => x"30c30c",
   14929 => x"30c30c",
   14930 => x"30c30c",
   14931 => x"30c30c",
   14932 => x"30c30c",
   14933 => x"30c30c",
   14934 => x"30c30c",
   14935 => x"30c30c",
   14936 => x"30c30c",
   14937 => x"30c30c",
   14938 => x"30c30c",
   14939 => x"30c30c",
   14940 => x"30c30c",
   14941 => x"30c30c",
   14942 => x"30c30c",
   14943 => x"30c30c",
   14944 => x"30c30c",
   14945 => x"30c30c",
   14946 => x"30c30c",
   14947 => x"30c30c",
   14948 => x"77ffff",
   14949 => x"ffffff",
   14950 => x"ffffff",
   14951 => x"ffffff",
   14952 => x"ffffff",
   14953 => x"ffffff",
   14954 => x"ffffff",
   14955 => x"ffffff",
   14956 => x"ffffff",
   14957 => x"ffffff",
   14958 => x"ffffff",
   14959 => x"ffffff",
   14960 => x"ffffff",
   14961 => x"ffffff",
   14962 => x"ffffff",
   14963 => x"ffffff",
   14964 => x"ffffff",
   14965 => x"ffffff",
   14966 => x"ffffff",
   14967 => x"ffffff",
   14968 => x"fea56a",
   14969 => x"ffffff",
   14970 => x"ffffff",
   14971 => x"ffffff",
   14972 => x"ffffff",
   14973 => x"ffffff",
   14974 => x"ffffff",
   14975 => x"ffffff",
   14976 => x"ffffff",
   14977 => x"ffffff",
   14978 => x"ffffff",
   14979 => x"ffffff",
   14980 => x"ffffff",
   14981 => x"ffffff",
   14982 => x"ffffff",
   14983 => x"ffffff",
   14984 => x"ffffff",
   14985 => x"ffffff",
   14986 => x"ffffff",
   14987 => x"ffffff",
   14988 => x"ffffff",
   14989 => x"ffffff",
   14990 => x"ffffff",
   14991 => x"ffffff",
   14992 => x"ffffff",
   14993 => x"ffffff",
   14994 => x"ffffff",
   14995 => x"ffffff",
   14996 => x"ffffff",
   14997 => x"ffffff",
   14998 => x"ffffff",
   14999 => x"ffffff",
   15000 => x"ffffff",
   15001 => x"ffffff",
   15002 => x"ffffff",
   15003 => x"ffffff",
   15004 => x"ffffff",
   15005 => x"ffffff",
   15006 => x"ffffff",
   15007 => x"ffffff",
   15008 => x"ffffff",
   15009 => x"ffffff",
   15010 => x"ffffff",
   15011 => x"ffffff",
   15012 => x"ffffff",
   15013 => x"ffffff",
   15014 => x"ffffff",
   15015 => x"ffffff",
   15016 => x"ffffff",
   15017 => x"ffffff",
   15018 => x"ffffff",
   15019 => x"ffffff",
   15020 => x"ffffff",
   15021 => x"ffffff",
   15022 => x"ffffff",
   15023 => x"ffffff",
   15024 => x"ffffff",
   15025 => x"ffffff",
   15026 => x"ffffff",
   15027 => x"ffffff",
   15028 => x"ffffff",
   15029 => x"ffffff",
   15030 => x"ffffff",
   15031 => x"ffffff",
   15032 => x"ffffff",
   15033 => x"ffffff",
   15034 => x"ffffff",
   15035 => x"ffffff",
   15036 => x"ffffff",
   15037 => x"ffffff",
   15038 => x"ffffff",
   15039 => x"ffffff",
   15040 => x"ffac30",
   15041 => x"c30c30",
   15042 => x"c30c30",
   15043 => x"c30c30",
   15044 => x"c30c30",
   15045 => x"c30c30",
   15046 => x"c30c30",
   15047 => x"c30c30",
   15048 => x"c30c30",
   15049 => x"c30c30",
   15050 => x"c30c30",
   15051 => x"c30c30",
   15052 => x"c30c30",
   15053 => x"c30c30",
   15054 => x"c30c30",
   15055 => x"c30c30",
   15056 => x"c30c30",
   15057 => x"c30c30",
   15058 => x"c30c30",
   15059 => x"c30c30",
   15060 => x"c30c30",
   15061 => x"c30c30",
   15062 => x"928f3c",
   15063 => x"f3cf3c",
   15064 => x"f3cf3c",
   15065 => x"f3cf3c",
   15066 => x"f3cf3c",
   15067 => x"f3cf3c",
   15068 => x"f3cf3c",
   15069 => x"f3cf3c",
   15070 => x"f3cf3c",
   15071 => x"f3cf3c",
   15072 => x"f3cf3c",
   15073 => x"f3cf3c",
   15074 => x"f3cf3c",
   15075 => x"f3cf3c",
   15076 => x"f3cf3c",
   15077 => x"f3cf3c",
   15078 => x"f3cf3c",
   15079 => x"f3cf3c",
   15080 => x"f3cf3c",
   15081 => x"f3cf3c",
   15082 => x"f3cf3c",
   15083 => x"f3cf3c",
   15084 => x"f3cf3c",
   15085 => x"f3cf3c",
   15086 => x"b0c30c",
   15087 => x"30c30c",
   15088 => x"30c30c",
   15089 => x"30c30c",
   15090 => x"30c30c",
   15091 => x"30c30c",
   15092 => x"30c30c",
   15093 => x"30c30c",
   15094 => x"30c30c",
   15095 => x"30c30c",
   15096 => x"30c30c",
   15097 => x"30c30c",
   15098 => x"30c30c",
   15099 => x"30c30c",
   15100 => x"30c30c",
   15101 => x"30c30c",
   15102 => x"30c30c",
   15103 => x"30c30c",
   15104 => x"30c30c",
   15105 => x"30c30c",
   15106 => x"30c30c",
   15107 => x"30c30c",
   15108 => x"77ffff",
   15109 => x"ffffff",
   15110 => x"ffffff",
   15111 => x"ffffff",
   15112 => x"ffffff",
   15113 => x"ffffff",
   15114 => x"ffffff",
   15115 => x"ffffff",
   15116 => x"ffffff",
   15117 => x"ffffff",
   15118 => x"ffffff",
   15119 => x"ffffff",
   15120 => x"ffffff",
   15121 => x"ffffff",
   15122 => x"ffffff",
   15123 => x"ffffff",
   15124 => x"ffffff",
   15125 => x"ffffff",
   15126 => x"ffffff",
   15127 => x"ffffff",
   15128 => x"a95abf",
   15129 => x"ffffff",
   15130 => x"ffffff",
   15131 => x"ffffff",
   15132 => x"ffffff",
   15133 => x"ffffff",
   15134 => x"ffffff",
   15135 => x"ffffff",
   15136 => x"ffffff",
   15137 => x"ffffff",
   15138 => x"ffffff",
   15139 => x"ffffff",
   15140 => x"ffffff",
   15141 => x"ffffff",
   15142 => x"ffffff",
   15143 => x"ffffff",
   15144 => x"ffffff",
   15145 => x"ffffff",
   15146 => x"ffffff",
   15147 => x"ffffff",
   15148 => x"ffffff",
   15149 => x"ffffff",
   15150 => x"ffffff",
   15151 => x"ffffff",
   15152 => x"ffffff",
   15153 => x"ffffff",
   15154 => x"ffffff",
   15155 => x"ffffff",
   15156 => x"ffffff",
   15157 => x"ffffff",
   15158 => x"ffffff",
   15159 => x"ffffff",
   15160 => x"ffffff",
   15161 => x"ffffff",
   15162 => x"ffffff",
   15163 => x"ffffff",
   15164 => x"ffffff",
   15165 => x"ffffff",
   15166 => x"ffffff",
   15167 => x"ffffff",
   15168 => x"ffffff",
   15169 => x"ffffff",
   15170 => x"ffffff",
   15171 => x"ffffff",
   15172 => x"ffffff",
   15173 => x"ffffff",
   15174 => x"ffffff",
   15175 => x"ffffff",
   15176 => x"ffffff",
   15177 => x"ffffff",
   15178 => x"ffffff",
   15179 => x"ffffff",
   15180 => x"ffffff",
   15181 => x"ffffff",
   15182 => x"ffffff",
   15183 => x"ffffff",
   15184 => x"ffffff",
   15185 => x"ffffff",
   15186 => x"ffffff",
   15187 => x"ffffff",
   15188 => x"ffffff",
   15189 => x"ffffff",
   15190 => x"ffffff",
   15191 => x"ffffff",
   15192 => x"ffffff",
   15193 => x"ffffff",
   15194 => x"ffffff",
   15195 => x"ffffff",
   15196 => x"ffffff",
   15197 => x"ffffff",
   15198 => x"ffffff",
   15199 => x"ffffff",
   15200 => x"ffac30",
   15201 => x"c30c30",
   15202 => x"c30c30",
   15203 => x"c30c30",
   15204 => x"c30c30",
   15205 => x"c30c30",
   15206 => x"c30c30",
   15207 => x"c30c30",
   15208 => x"c30c30",
   15209 => x"c30c30",
   15210 => x"c30c30",
   15211 => x"c30c30",
   15212 => x"c30c30",
   15213 => x"c30c30",
   15214 => x"c30c30",
   15215 => x"c30c30",
   15216 => x"c30c30",
   15217 => x"c30c30",
   15218 => x"c30c30",
   15219 => x"c30c30",
   15220 => x"c30c30",
   15221 => x"c30c30",
   15222 => x"928f3c",
   15223 => x"f3cf3c",
   15224 => x"f3cf3c",
   15225 => x"f3cf3c",
   15226 => x"f3cf3c",
   15227 => x"f3cf3c",
   15228 => x"f3cf3c",
   15229 => x"f3cf3c",
   15230 => x"f3cf3c",
   15231 => x"f3cf3c",
   15232 => x"f3cf3c",
   15233 => x"f3cf3c",
   15234 => x"f3cf3c",
   15235 => x"f3cf3c",
   15236 => x"f3cf3c",
   15237 => x"f3cf3c",
   15238 => x"f3cf3c",
   15239 => x"f3cf3c",
   15240 => x"f3cf3c",
   15241 => x"f3cf3c",
   15242 => x"f3cf3c",
   15243 => x"f3cf3c",
   15244 => x"f3cf3c",
   15245 => x"f3cf3c",
   15246 => x"b0c30c",
   15247 => x"30c30c",
   15248 => x"30c30c",
   15249 => x"30c30c",
   15250 => x"30c30c",
   15251 => x"30c30c",
   15252 => x"30c30c",
   15253 => x"30c30c",
   15254 => x"30c30c",
   15255 => x"30c30c",
   15256 => x"30c30c",
   15257 => x"30c30c",
   15258 => x"30c30c",
   15259 => x"30c30c",
   15260 => x"30c30c",
   15261 => x"30c30c",
   15262 => x"30c30c",
   15263 => x"30c30c",
   15264 => x"30c30c",
   15265 => x"30c30c",
   15266 => x"30c30c",
   15267 => x"30c30c",
   15268 => x"77ffff",
   15269 => x"ffffff",
   15270 => x"ffffff",
   15271 => x"ffffff",
   15272 => x"ffffff",
   15273 => x"ffffff",
   15274 => x"ffffff",
   15275 => x"ffffff",
   15276 => x"ffffff",
   15277 => x"ffffff",
   15278 => x"ffffff",
   15279 => x"ffffff",
   15280 => x"ffffff",
   15281 => x"ffffff",
   15282 => x"ffffff",
   15283 => x"ffffff",
   15284 => x"ffffff",
   15285 => x"ffffff",
   15286 => x"ffffff",
   15287 => x"ffffea",
   15288 => x"56afff",
   15289 => x"ffffff",
   15290 => x"ffffff",
   15291 => x"ffffff",
   15292 => x"ffffff",
   15293 => x"ffffff",
   15294 => x"ffffff",
   15295 => x"ffffff",
   15296 => x"ffffff",
   15297 => x"ffffff",
   15298 => x"ffffff",
   15299 => x"ffffff",
   15300 => x"ffffff",
   15301 => x"ffffff",
   15302 => x"ffffff",
   15303 => x"ffffff",
   15304 => x"ffffff",
   15305 => x"ffffff",
   15306 => x"ffffff",
   15307 => x"ffffff",
   15308 => x"ffffff",
   15309 => x"ffffff",
   15310 => x"ffffff",
   15311 => x"ffffff",
   15312 => x"ffffff",
   15313 => x"ffffff",
   15314 => x"ffffff",
   15315 => x"ffffff",
   15316 => x"ffffff",
   15317 => x"ffffff",
   15318 => x"ffffff",
   15319 => x"ffffff",
   15320 => x"ffffff",
   15321 => x"ffffff",
   15322 => x"ffffff",
   15323 => x"ffffff",
   15324 => x"ffffff",
   15325 => x"ffffff",
   15326 => x"ffffff",
   15327 => x"ffffff",
   15328 => x"ffffff",
   15329 => x"ffffff",
   15330 => x"ffffff",
   15331 => x"ffffff",
   15332 => x"ffffff",
   15333 => x"ffffff",
   15334 => x"ffffff",
   15335 => x"ffffff",
   15336 => x"ffffff",
   15337 => x"ffffff",
   15338 => x"ffffff",
   15339 => x"ffffff",
   15340 => x"ffffff",
   15341 => x"ffffff",
   15342 => x"ffffff",
   15343 => x"ffffff",
   15344 => x"ffffff",
   15345 => x"ffffff",
   15346 => x"ffffff",
   15347 => x"ffffff",
   15348 => x"ffffff",
   15349 => x"ffffff",
   15350 => x"ffffff",
   15351 => x"ffffff",
   15352 => x"ffffff",
   15353 => x"ffffff",
   15354 => x"ffffff",
   15355 => x"ffffff",
   15356 => x"ffffff",
   15357 => x"ffffff",
   15358 => x"ffffff",
   15359 => x"ffffff",
   15360 => x"ffac30",
   15361 => x"c30c30",
   15362 => x"c30c30",
   15363 => x"c30c30",
   15364 => x"c30c30",
   15365 => x"c30c30",
   15366 => x"c30c30",
   15367 => x"c30c30",
   15368 => x"c30c30",
   15369 => x"c30c30",
   15370 => x"c30c30",
   15371 => x"c30c30",
   15372 => x"c30c30",
   15373 => x"c30c30",
   15374 => x"c30c30",
   15375 => x"c30c30",
   15376 => x"c30c30",
   15377 => x"c30c30",
   15378 => x"c30c30",
   15379 => x"c30c30",
   15380 => x"c30c30",
   15381 => x"c30c30",
   15382 => x"928f3c",
   15383 => x"f3cf3c",
   15384 => x"f3cf3c",
   15385 => x"f3cf3c",
   15386 => x"f3cf3c",
   15387 => x"f3cf3c",
   15388 => x"f3cf3c",
   15389 => x"f3cf3c",
   15390 => x"f3cf3c",
   15391 => x"f3cf3c",
   15392 => x"f3cf3c",
   15393 => x"f3cf3c",
   15394 => x"f3cf3c",
   15395 => x"f3cf3c",
   15396 => x"f3cf3c",
   15397 => x"f3cf3c",
   15398 => x"f3cf3c",
   15399 => x"f3cf3c",
   15400 => x"f3cf3c",
   15401 => x"f3cf3c",
   15402 => x"f3cf3c",
   15403 => x"f3cf3c",
   15404 => x"f3cf3c",
   15405 => x"f3cf3c",
   15406 => x"f0c30c",
   15407 => x"30c30c",
   15408 => x"30c30c",
   15409 => x"30c30c",
   15410 => x"30c30c",
   15411 => x"30c30c",
   15412 => x"30c30c",
   15413 => x"30c30c",
   15414 => x"30c30c",
   15415 => x"30c30c",
   15416 => x"30c30c",
   15417 => x"30c30c",
   15418 => x"30c30c",
   15419 => x"30c30c",
   15420 => x"30c30c",
   15421 => x"30c30c",
   15422 => x"30c30c",
   15423 => x"30c30c",
   15424 => x"30c30c",
   15425 => x"30c30c",
   15426 => x"30c30c",
   15427 => x"30c30c",
   15428 => x"77ffff",
   15429 => x"ffffff",
   15430 => x"ffffff",
   15431 => x"ffffff",
   15432 => x"ffffff",
   15433 => x"ffffff",
   15434 => x"ffffff",
   15435 => x"ffffff",
   15436 => x"ffffff",
   15437 => x"ffffff",
   15438 => x"ffffff",
   15439 => x"ffffff",
   15440 => x"ffffff",
   15441 => x"ffffff",
   15442 => x"ffffff",
   15443 => x"ffffff",
   15444 => x"ffffff",
   15445 => x"ffffff",
   15446 => x"ffffff",
   15447 => x"fffa95",
   15448 => x"abffff",
   15449 => x"ffffff",
   15450 => x"ffffff",
   15451 => x"ffffff",
   15452 => x"ffffff",
   15453 => x"ffffff",
   15454 => x"ffffff",
   15455 => x"ffffff",
   15456 => x"ffffff",
   15457 => x"ffffff",
   15458 => x"ffffff",
   15459 => x"ffffff",
   15460 => x"ffffff",
   15461 => x"ffffff",
   15462 => x"ffffff",
   15463 => x"ffffff",
   15464 => x"ffffff",
   15465 => x"ffffff",
   15466 => x"ffffff",
   15467 => x"ffffff",
   15468 => x"ffffff",
   15469 => x"ffffff",
   15470 => x"ffffff",
   15471 => x"ffffff",
   15472 => x"ffffff",
   15473 => x"ffffff",
   15474 => x"ffffff",
   15475 => x"ffffff",
   15476 => x"ffffff",
   15477 => x"ffffff",
   15478 => x"ffffff",
   15479 => x"ffffff",
   15480 => x"ffffff",
   15481 => x"ffffff",
   15482 => x"ffffff",
   15483 => x"ffffff",
   15484 => x"ffffff",
   15485 => x"ffffff",
   15486 => x"ffffff",
   15487 => x"ffffff",
   15488 => x"ffffff",
   15489 => x"ffffff",
   15490 => x"ffffff",
   15491 => x"ffffff",
   15492 => x"ffffff",
   15493 => x"ffffff",
   15494 => x"ffffff",
   15495 => x"ffffff",
   15496 => x"ffffff",
   15497 => x"ffffff",
   15498 => x"ffffff",
   15499 => x"ffffff",
   15500 => x"ffffff",
   15501 => x"ffffff",
   15502 => x"ffffff",
   15503 => x"ffffff",
   15504 => x"ffffff",
   15505 => x"ffffff",
   15506 => x"ffffff",
   15507 => x"ffffff",
   15508 => x"ffffff",
   15509 => x"ffffff",
   15510 => x"ffffff",
   15511 => x"ffffff",
   15512 => x"ffffff",
   15513 => x"ffffff",
   15514 => x"ffffff",
   15515 => x"ffffff",
   15516 => x"ffffff",
   15517 => x"ffffff",
   15518 => x"ffffff",
   15519 => x"ffffff",
   15520 => x"ffac30",
   15521 => x"c30c30",
   15522 => x"c30c30",
   15523 => x"c30c30",
   15524 => x"c30c30",
   15525 => x"c30c30",
   15526 => x"c30c30",
   15527 => x"c30c30",
   15528 => x"c30c30",
   15529 => x"c30c30",
   15530 => x"c30c30",
   15531 => x"c30c30",
   15532 => x"c30c30",
   15533 => x"c30c30",
   15534 => x"c30c30",
   15535 => x"c30c30",
   15536 => x"c30c30",
   15537 => x"c30c30",
   15538 => x"c30c30",
   15539 => x"c30c30",
   15540 => x"c30c30",
   15541 => x"c30c30",
   15542 => x"92cf3c",
   15543 => x"f3cf3c",
   15544 => x"f3cf3c",
   15545 => x"f3cf3c",
   15546 => x"f3cf3c",
   15547 => x"f3cf3c",
   15548 => x"f3cf3c",
   15549 => x"f3cf3c",
   15550 => x"f3cf3c",
   15551 => x"f3cf3c",
   15552 => x"f3cf3c",
   15553 => x"f3cf3c",
   15554 => x"f3cf3c",
   15555 => x"f3cf3c",
   15556 => x"f3cf3c",
   15557 => x"f3cf3c",
   15558 => x"f3cf3c",
   15559 => x"f3cf3c",
   15560 => x"f3cf3c",
   15561 => x"f3cf3c",
   15562 => x"f3cf3c",
   15563 => x"f3cf3c",
   15564 => x"f3cf3c",
   15565 => x"f3cf3c",
   15566 => x"f0c30c",
   15567 => x"30c30c",
   15568 => x"30c30c",
   15569 => x"30c30c",
   15570 => x"30c30c",
   15571 => x"30c30c",
   15572 => x"30c30c",
   15573 => x"30c30c",
   15574 => x"30c30c",
   15575 => x"30c30c",
   15576 => x"30c30c",
   15577 => x"30c30c",
   15578 => x"30c30c",
   15579 => x"30c30c",
   15580 => x"30c30c",
   15581 => x"30c30c",
   15582 => x"30c30c",
   15583 => x"30c30c",
   15584 => x"30c30c",
   15585 => x"30c30c",
   15586 => x"30c30c",
   15587 => x"30c30c",
   15588 => x"76efff",
   15589 => x"ffffff",
   15590 => x"ffffff",
   15591 => x"ffffff",
   15592 => x"ffffff",
   15593 => x"ffffff",
   15594 => x"ffffff",
   15595 => x"ffffff",
   15596 => x"ffffff",
   15597 => x"ffffff",
   15598 => x"ffffff",
   15599 => x"ffffff",
   15600 => x"ffffff",
   15601 => x"ffffff",
   15602 => x"ffffff",
   15603 => x"ffffff",
   15604 => x"ffffff",
   15605 => x"ffffff",
   15606 => x"ffffff",
   15607 => x"fea56a",
   15608 => x"ffffff",
   15609 => x"ffffff",
   15610 => x"ffffff",
   15611 => x"ffffff",
   15612 => x"ffffff",
   15613 => x"ffffff",
   15614 => x"ffffff",
   15615 => x"ffffff",
   15616 => x"ffffff",
   15617 => x"ffffff",
   15618 => x"ffffff",
   15619 => x"ffffff",
   15620 => x"ffffff",
   15621 => x"ffffff",
   15622 => x"ffffff",
   15623 => x"ffffff",
   15624 => x"ffffff",
   15625 => x"ffffff",
   15626 => x"ffffff",
   15627 => x"ffffff",
   15628 => x"ffffff",
   15629 => x"ffffff",
   15630 => x"ffffff",
   15631 => x"ffffff",
   15632 => x"ffffff",
   15633 => x"ffffff",
   15634 => x"ffffff",
   15635 => x"ffffff",
   15636 => x"ffffff",
   15637 => x"ffffff",
   15638 => x"ffffff",
   15639 => x"ffffff",
   15640 => x"ffffff",
   15641 => x"ffffff",
   15642 => x"ffffff",
   15643 => x"ffffff",
   15644 => x"ffffff",
   15645 => x"ffffff",
   15646 => x"ffffff",
   15647 => x"ffffff",
   15648 => x"ffffff",
   15649 => x"ffffff",
   15650 => x"ffffff",
   15651 => x"ffffff",
   15652 => x"ffffff",
   15653 => x"ffffff",
   15654 => x"ffffff",
   15655 => x"ffffff",
   15656 => x"ffffff",
   15657 => x"ffffff",
   15658 => x"ffffff",
   15659 => x"ffffff",
   15660 => x"ffffff",
   15661 => x"ffffff",
   15662 => x"ffffff",
   15663 => x"ffffff",
   15664 => x"ffffff",
   15665 => x"ffffff",
   15666 => x"ffffff",
   15667 => x"ffffff",
   15668 => x"ffffff",
   15669 => x"ffffff",
   15670 => x"ffffff",
   15671 => x"ffffff",
   15672 => x"ffffff",
   15673 => x"ffffff",
   15674 => x"ffffff",
   15675 => x"ffffff",
   15676 => x"ffffff",
   15677 => x"ffffff",
   15678 => x"ffffff",
   15679 => x"ffffff",
   15680 => x"ffac30",
   15681 => x"c30c30",
   15682 => x"c30c30",
   15683 => x"c30c30",
   15684 => x"c30c30",
   15685 => x"c30c30",
   15686 => x"c30c30",
   15687 => x"c30c30",
   15688 => x"c30c30",
   15689 => x"c30c30",
   15690 => x"c30c30",
   15691 => x"c30c30",
   15692 => x"c30c30",
   15693 => x"c30c30",
   15694 => x"c30c30",
   15695 => x"c30c30",
   15696 => x"c30c30",
   15697 => x"c30c30",
   15698 => x"c30c30",
   15699 => x"c30c30",
   15700 => x"c30c30",
   15701 => x"c30c30",
   15702 => x"92cf3c",
   15703 => x"f3cf3c",
   15704 => x"f3cf3c",
   15705 => x"f3cf3c",
   15706 => x"f3cf3c",
   15707 => x"f3cf3c",
   15708 => x"f3cf3c",
   15709 => x"f3cf3c",
   15710 => x"f3cf3c",
   15711 => x"f3cf3c",
   15712 => x"f3cf3c",
   15713 => x"f3cf3c",
   15714 => x"f3cf3c",
   15715 => x"f3cf3c",
   15716 => x"f3cf3c",
   15717 => x"f3cf3c",
   15718 => x"f3cf3c",
   15719 => x"f3cf3c",
   15720 => x"f3cf3c",
   15721 => x"f3cf3c",
   15722 => x"f3cf3c",
   15723 => x"f3cf3c",
   15724 => x"f3cf3c",
   15725 => x"f3cf3c",
   15726 => x"f1c30c",
   15727 => x"30c30c",
   15728 => x"30c30c",
   15729 => x"30c30c",
   15730 => x"30c30c",
   15731 => x"30c30c",
   15732 => x"30c30c",
   15733 => x"30c30c",
   15734 => x"30c30c",
   15735 => x"30c30c",
   15736 => x"30c30c",
   15737 => x"30c30c",
   15738 => x"30c30c",
   15739 => x"30c30c",
   15740 => x"30c30c",
   15741 => x"30c30c",
   15742 => x"30c30c",
   15743 => x"30c30c",
   15744 => x"30c30c",
   15745 => x"30c30c",
   15746 => x"30c30c",
   15747 => x"30c30c",
   15748 => x"32efff",
   15749 => x"ffffff",
   15750 => x"ffffff",
   15751 => x"ffffff",
   15752 => x"ffffff",
   15753 => x"ffffff",
   15754 => x"ffffff",
   15755 => x"ffffff",
   15756 => x"ffffff",
   15757 => x"ffffff",
   15758 => x"ffffff",
   15759 => x"ffffff",
   15760 => x"ffffff",
   15761 => x"ffffff",
   15762 => x"ffffff",
   15763 => x"ffffff",
   15764 => x"ffffff",
   15765 => x"ffffff",
   15766 => x"ffffff",
   15767 => x"a95abf",
   15768 => x"ffffff",
   15769 => x"ffffff",
   15770 => x"ffffff",
   15771 => x"ffffff",
   15772 => x"ffffff",
   15773 => x"ffffff",
   15774 => x"ffffff",
   15775 => x"ffffff",
   15776 => x"ffffff",
   15777 => x"ffffff",
   15778 => x"ffffff",
   15779 => x"ffffff",
   15780 => x"ffffff",
   15781 => x"ffffff",
   15782 => x"ffffff",
   15783 => x"ffffff",
   15784 => x"ffffff",
   15785 => x"ffffff",
   15786 => x"ffffff",
   15787 => x"ffffff",
   15788 => x"ffffff",
   15789 => x"ffffff",
   15790 => x"ffffff",
   15791 => x"ffffff",
   15792 => x"ffffff",
   15793 => x"ffffff",
   15794 => x"ffffff",
   15795 => x"ffffff",
   15796 => x"ffffff",
   15797 => x"ffffff",
   15798 => x"ffffff",
   15799 => x"ffffff",
   15800 => x"ffffff",
   15801 => x"ffffff",
   15802 => x"ffffff",
   15803 => x"ffffff",
   15804 => x"ffffff",
   15805 => x"ffffff",
   15806 => x"ffffff",
   15807 => x"ffffff",
   15808 => x"ffffff",
   15809 => x"ffffff",
   15810 => x"ffffff",
   15811 => x"ffffff",
   15812 => x"ffffff",
   15813 => x"ffffff",
   15814 => x"ffffff",
   15815 => x"ffffff",
   15816 => x"ffffff",
   15817 => x"ffffff",
   15818 => x"ffffff",
   15819 => x"ffffff",
   15820 => x"ffffff",
   15821 => x"ffffff",
   15822 => x"ffffff",
   15823 => x"ffffff",
   15824 => x"ffffff",
   15825 => x"ffffff",
   15826 => x"ffffff",
   15827 => x"ffffff",
   15828 => x"ffffff",
   15829 => x"ffffff",
   15830 => x"ffffff",
   15831 => x"ffffff",
   15832 => x"ffffff",
   15833 => x"ffffff",
   15834 => x"ffffff",
   15835 => x"ffffff",
   15836 => x"ffffff",
   15837 => x"ffffff",
   15838 => x"ffffff",
   15839 => x"ffffff",
   15840 => x"ffac30",
   15841 => x"c30c30",
   15842 => x"c30c30",
   15843 => x"c30c30",
   15844 => x"c30c30",
   15845 => x"c30c30",
   15846 => x"c30c30",
   15847 => x"c30c30",
   15848 => x"c30c30",
   15849 => x"c30c30",
   15850 => x"c30c30",
   15851 => x"c30c30",
   15852 => x"c30c30",
   15853 => x"c30c30",
   15854 => x"c30c30",
   15855 => x"c30c30",
   15856 => x"c30c30",
   15857 => x"c30c30",
   15858 => x"c30c30",
   15859 => x"c30c30",
   15860 => x"c30c30",
   15861 => x"c30c30",
   15862 => x"92cf3c",
   15863 => x"f3cf3c",
   15864 => x"f3cf3c",
   15865 => x"f3cf3c",
   15866 => x"f3cf3c",
   15867 => x"f3cf3c",
   15868 => x"f3cf3c",
   15869 => x"f3cf3c",
   15870 => x"f3cf3c",
   15871 => x"f3cf3c",
   15872 => x"f3cb2c",
   15873 => x"b2cb2c",
   15874 => x"b2cb2c",
   15875 => x"b2cb2c",
   15876 => x"b3cf3c",
   15877 => x"f3cf3c",
   15878 => x"f3cf3c",
   15879 => x"f3cf3c",
   15880 => x"f3cf3c",
   15881 => x"f3cf3c",
   15882 => x"f3cf3c",
   15883 => x"f3cf3c",
   15884 => x"f3cf3c",
   15885 => x"f3cf3c",
   15886 => x"f1c30c",
   15887 => x"30c30c",
   15888 => x"30c30c",
   15889 => x"30c30c",
   15890 => x"30c30c",
   15891 => x"30c30c",
   15892 => x"30c30c",
   15893 => x"30c30c",
   15894 => x"30c30c",
   15895 => x"30c30c",
   15896 => x"30c30c",
   15897 => x"30c30c",
   15898 => x"30c30c",
   15899 => x"30c30c",
   15900 => x"30c30c",
   15901 => x"30c30c",
   15902 => x"30c30c",
   15903 => x"30c30c",
   15904 => x"30c30c",
   15905 => x"30c30c",
   15906 => x"30c30c",
   15907 => x"30c30c",
   15908 => x"32efff",
   15909 => x"ffffff",
   15910 => x"ffffff",
   15911 => x"ffffff",
   15912 => x"ffffff",
   15913 => x"ffffff",
   15914 => x"ffffff",
   15915 => x"ffffff",
   15916 => x"ffffff",
   15917 => x"ffffff",
   15918 => x"ffffff",
   15919 => x"ffffff",
   15920 => x"ffffff",
   15921 => x"ffffff",
   15922 => x"ffffff",
   15923 => x"ffffff",
   15924 => x"ffffff",
   15925 => x"ffffff",
   15926 => x"ffffea",
   15927 => x"56afff",
   15928 => x"ffffff",
   15929 => x"ffffff",
   15930 => x"ffffff",
   15931 => x"ffffff",
   15932 => x"ffffff",
   15933 => x"ffffff",
   15934 => x"ffffff",
   15935 => x"ffffff",
   15936 => x"ffffff",
   15937 => x"ffffff",
   15938 => x"ffffff",
   15939 => x"ffffff",
   15940 => x"ffffff",
   15941 => x"ffffff",
   15942 => x"ffffff",
   15943 => x"ffffff",
   15944 => x"ffffff",
   15945 => x"ffffff",
   15946 => x"ffffff",
   15947 => x"ffffff",
   15948 => x"ffffff",
   15949 => x"ffffff",
   15950 => x"ffffff",
   15951 => x"ffffff",
   15952 => x"ffffff",
   15953 => x"ffffff",
   15954 => x"ffffff",
   15955 => x"ffffff",
   15956 => x"ffffff",
   15957 => x"ffffff",
   15958 => x"ffffff",
   15959 => x"ffffff",
   15960 => x"ffffff",
   15961 => x"ffffff",
   15962 => x"ffffff",
   15963 => x"ffffff",
   15964 => x"ffffff",
   15965 => x"ffffff",
   15966 => x"ffffff",
   15967 => x"ffffff",
   15968 => x"ffffff",
   15969 => x"ffffff",
   15970 => x"ffffff",
   15971 => x"ffffff",
   15972 => x"ffffff",
   15973 => x"ffffff",
   15974 => x"ffffff",
   15975 => x"ffffff",
   15976 => x"ffffff",
   15977 => x"ffffff",
   15978 => x"ffffff",
   15979 => x"ffffff",
   15980 => x"ffffff",
   15981 => x"ffffff",
   15982 => x"ffffff",
   15983 => x"ffffff",
   15984 => x"ffffff",
   15985 => x"ffffff",
   15986 => x"ffffff",
   15987 => x"ffffff",
   15988 => x"ffffff",
   15989 => x"ffffff",
   15990 => x"ffffff",
   15991 => x"ffffff",
   15992 => x"ffffff",
   15993 => x"ffffff",
   15994 => x"ffffff",
   15995 => x"ffffff",
   15996 => x"ffffff",
   15997 => x"ffffff",
   15998 => x"ffffff",
   15999 => x"ffffff",
   16000 => x"ff5c30",
   16001 => x"c30c30",
   16002 => x"c30c30",
   16003 => x"c30c30",
   16004 => x"c30c30",
   16005 => x"c30c30",
   16006 => x"c30c30",
   16007 => x"c30c30",
   16008 => x"c30c30",
   16009 => x"c30c30",
   16010 => x"c30c30",
   16011 => x"c30c30",
   16012 => x"c30c30",
   16013 => x"c30c30",
   16014 => x"c30c30",
   16015 => x"c30c30",
   16016 => x"c30c30",
   16017 => x"c30c30",
   16018 => x"c30c30",
   16019 => x"c30c30",
   16020 => x"c30c30",
   16021 => x"c30c30",
   16022 => x"92cf3c",
   16023 => x"f3cf3c",
   16024 => x"f3cf3c",
   16025 => x"f3cf3c",
   16026 => x"f3cf3c",
   16027 => x"f3cf3c",
   16028 => x"f3cf3c",
   16029 => x"f3cf3c",
   16030 => x"f3cb2c",
   16031 => x"b6d75d",
   16032 => x"7aebae",
   16033 => x"baebae",
   16034 => x"baebae",
   16035 => x"baebae",
   16036 => x"bae75d",
   16037 => x"75d76c",
   16038 => x"b3cf3c",
   16039 => x"f3cf3c",
   16040 => x"f3cf3c",
   16041 => x"f3cf3c",
   16042 => x"f3cf3c",
   16043 => x"f3cf3c",
   16044 => x"f3cf3c",
   16045 => x"f3cf3c",
   16046 => x"f1c30c",
   16047 => x"30c30c",
   16048 => x"30c30c",
   16049 => x"30c30c",
   16050 => x"30c30c",
   16051 => x"30c30c",
   16052 => x"30c30c",
   16053 => x"30c30c",
   16054 => x"30c30c",
   16055 => x"30c30c",
   16056 => x"30c30c",
   16057 => x"30c30c",
   16058 => x"30c30c",
   16059 => x"30c30c",
   16060 => x"30c30c",
   16061 => x"30c30c",
   16062 => x"30c30c",
   16063 => x"30c30c",
   16064 => x"30c30c",
   16065 => x"30c30c",
   16066 => x"30c30c",
   16067 => x"30c30c",
   16068 => x"32efff",
   16069 => x"ffffff",
   16070 => x"ffffff",
   16071 => x"ffffff",
   16072 => x"ffffff",
   16073 => x"ffffff",
   16074 => x"ffffff",
   16075 => x"ffffff",
   16076 => x"ffffff",
   16077 => x"ffffff",
   16078 => x"ffffff",
   16079 => x"ffffff",
   16080 => x"ffffff",
   16081 => x"ffffff",
   16082 => x"ffffff",
   16083 => x"ffffff",
   16084 => x"ffffff",
   16085 => x"ffffff",
   16086 => x"fffa95",
   16087 => x"abffff",
   16088 => x"ffffff",
   16089 => x"ffffff",
   16090 => x"ffffff",
   16091 => x"ffffff",
   16092 => x"ffffff",
   16093 => x"ffffff",
   16094 => x"ffffff",
   16095 => x"ffffff",
   16096 => x"ffffff",
   16097 => x"ffffff",
   16098 => x"ffffff",
   16099 => x"ffffff",
   16100 => x"ffffff",
   16101 => x"ffffff",
   16102 => x"ffffff",
   16103 => x"ffffff",
   16104 => x"ffffff",
   16105 => x"ffffff",
   16106 => x"ffffff",
   16107 => x"ffffff",
   16108 => x"ffffff",
   16109 => x"ffffff",
   16110 => x"ffffff",
   16111 => x"ffffff",
   16112 => x"ffffff",
   16113 => x"ffffff",
   16114 => x"ffffff",
   16115 => x"ffffff",
   16116 => x"ffffff",
   16117 => x"ffffff",
   16118 => x"ffffff",
   16119 => x"ffffff",
   16120 => x"ffffff",
   16121 => x"ffffff",
   16122 => x"ffffff",
   16123 => x"ffffff",
   16124 => x"ffffff",
   16125 => x"ffffff",
   16126 => x"ffffff",
   16127 => x"ffffff",
   16128 => x"ffffff",
   16129 => x"ffffff",
   16130 => x"ffffff",
   16131 => x"ffffff",
   16132 => x"ffffff",
   16133 => x"ffffff",
   16134 => x"ffffff",
   16135 => x"ffffff",
   16136 => x"ffffff",
   16137 => x"ffffff",
   16138 => x"ffffff",
   16139 => x"ffffff",
   16140 => x"ffffff",
   16141 => x"ffffff",
   16142 => x"ffffff",
   16143 => x"ffffff",
   16144 => x"ffffff",
   16145 => x"ffffff",
   16146 => x"ffffff",
   16147 => x"ffffff",
   16148 => x"ffffff",
   16149 => x"ffffff",
   16150 => x"ffffff",
   16151 => x"ffffff",
   16152 => x"ffffff",
   16153 => x"ffffff",
   16154 => x"ffffff",
   16155 => x"ffffff",
   16156 => x"ffffff",
   16157 => x"ffffff",
   16158 => x"ffffff",
   16159 => x"ffffff",
   16160 => x"ff5c30",
   16161 => x"c30c30",
   16162 => x"c30c30",
   16163 => x"c30c30",
   16164 => x"c30c30",
   16165 => x"c30c30",
   16166 => x"c30c30",
   16167 => x"c30c30",
   16168 => x"c30c30",
   16169 => x"c30c30",
   16170 => x"c30c30",
   16171 => x"c30c30",
   16172 => x"c30c30",
   16173 => x"c30c30",
   16174 => x"c30c30",
   16175 => x"c30c30",
   16176 => x"c30c30",
   16177 => x"c30c30",
   16178 => x"c30c30",
   16179 => x"c30c30",
   16180 => x"c30c30",
   16181 => x"c30c30",
   16182 => x"92cf3c",
   16183 => x"f3cf3c",
   16184 => x"f3cf3c",
   16185 => x"f3cf3c",
   16186 => x"f3cf3c",
   16187 => x"f3cf3c",
   16188 => x"f3cf3c",
   16189 => x"b2cb6d",
   16190 => x"b6ebbf",
   16191 => x"ffffff",
   16192 => x"ffffff",
   16193 => x"ffffff",
   16194 => x"ffffff",
   16195 => x"ffffff",
   16196 => x"ffffff",
   16197 => x"ffffff",
   16198 => x"bae75d",
   16199 => x"b2cb3c",
   16200 => x"f3cf3c",
   16201 => x"f3cf3c",
   16202 => x"f3cf3c",
   16203 => x"f3cf3c",
   16204 => x"f3cf3c",
   16205 => x"f3cf3c",
   16206 => x"f1c30c",
   16207 => x"30c30c",
   16208 => x"30c30c",
   16209 => x"30c30c",
   16210 => x"30c30c",
   16211 => x"30c30c",
   16212 => x"30c30c",
   16213 => x"30c30c",
   16214 => x"30c30c",
   16215 => x"30c30c",
   16216 => x"30c30c",
   16217 => x"30c30c",
   16218 => x"30c30c",
   16219 => x"30c30c",
   16220 => x"30c30c",
   16221 => x"30c30c",
   16222 => x"30c30c",
   16223 => x"30c30c",
   16224 => x"30c30c",
   16225 => x"30c30c",
   16226 => x"30c30c",
   16227 => x"30c30c",
   16228 => x"32efff",
   16229 => x"ffffff",
   16230 => x"ffffff",
   16231 => x"ffffff",
   16232 => x"ffffff",
   16233 => x"ffffff",
   16234 => x"ffffff",
   16235 => x"ffffff",
   16236 => x"ffffff",
   16237 => x"ffffff",
   16238 => x"ffffff",
   16239 => x"ffffff",
   16240 => x"ffffff",
   16241 => x"ffffff",
   16242 => x"ffffff",
   16243 => x"ffffff",
   16244 => x"ffffff",
   16245 => x"ffffff",
   16246 => x"fea56a",
   16247 => x"ffffff",
   16248 => x"ffffff",
   16249 => x"ffffff",
   16250 => x"ffffff",
   16251 => x"ffffff",
   16252 => x"ffffff",
   16253 => x"ffffff",
   16254 => x"ffffff",
   16255 => x"ffffff",
   16256 => x"ffffff",
   16257 => x"ffffff",
   16258 => x"ffffff",
   16259 => x"ffffff",
   16260 => x"ffffff",
   16261 => x"ffffff",
   16262 => x"ffffff",
   16263 => x"ffffff",
   16264 => x"ffffff",
   16265 => x"ffffff",
   16266 => x"ffffff",
   16267 => x"ffffff",
   16268 => x"ffffff",
   16269 => x"ffffff",
   16270 => x"ffffff",
   16271 => x"ffffff",
   16272 => x"ffffff",
   16273 => x"ffffff",
   16274 => x"ffffff",
   16275 => x"ffffff",
   16276 => x"ffffff",
   16277 => x"ffffff",
   16278 => x"ffffff",
   16279 => x"ffffff",
   16280 => x"ffffff",
   16281 => x"ffffff",
   16282 => x"ffffff",
   16283 => x"ffffff",
   16284 => x"ffffff",
   16285 => x"ffffff",
   16286 => x"ffffff",
   16287 => x"ffffff",
   16288 => x"ffffff",
   16289 => x"ffffff",
   16290 => x"ffffff",
   16291 => x"ffffff",
   16292 => x"ffffff",
   16293 => x"ffffff",
   16294 => x"ffffff",
   16295 => x"ffffff",
   16296 => x"ffffff",
   16297 => x"ffffff",
   16298 => x"ffffff",
   16299 => x"ffffff",
   16300 => x"ffffff",
   16301 => x"ffffff",
   16302 => x"ffffff",
   16303 => x"ffffff",
   16304 => x"ffffff",
   16305 => x"ffffff",
   16306 => x"ffffff",
   16307 => x"ffffff",
   16308 => x"ffffff",
   16309 => x"ffffff",
   16310 => x"ffffff",
   16311 => x"ffffff",
   16312 => x"ffffff",
   16313 => x"ffffff",
   16314 => x"ffffff",
   16315 => x"ffffff",
   16316 => x"ffffff",
   16317 => x"ffffff",
   16318 => x"ffffff",
   16319 => x"ffffff",
   16320 => x"ff5c30",
   16321 => x"c30c30",
   16322 => x"c30c30",
   16323 => x"c30c30",
   16324 => x"c30c30",
   16325 => x"c30c30",
   16326 => x"c30c30",
   16327 => x"c30c30",
   16328 => x"c30c30",
   16329 => x"c30c30",
   16330 => x"c30c30",
   16331 => x"c30c30",
   16332 => x"c30c30",
   16333 => x"c30c30",
   16334 => x"c30c30",
   16335 => x"c30c30",
   16336 => x"c30c30",
   16337 => x"c30c30",
   16338 => x"c30c30",
   16339 => x"c30c30",
   16340 => x"c30c30",
   16341 => x"c30c30",
   16342 => x"a2cf3c",
   16343 => x"f3cf3c",
   16344 => x"f3cf3c",
   16345 => x"f3cf3c",
   16346 => x"f3cf3c",
   16347 => x"f3cf3c",
   16348 => x"f2c76d",
   16349 => x"bbffff",
   16350 => x"ffffff",
   16351 => x"ffffff",
   16352 => x"ffffff",
   16353 => x"ffffff",
   16354 => x"ffffff",
   16355 => x"ffffff",
   16356 => x"ffffff",
   16357 => x"ffffff",
   16358 => x"ffffff",
   16359 => x"feeb9d",
   16360 => x"76cb3c",
   16361 => x"f3cf3c",
   16362 => x"f3cf3c",
   16363 => x"f3cf3c",
   16364 => x"f3cf3c",
   16365 => x"f3cf3c",
   16366 => x"f2c30c",
   16367 => x"30c30c",
   16368 => x"30c30c",
   16369 => x"30c30c",
   16370 => x"30c30c",
   16371 => x"30c30c",
   16372 => x"30c30c",
   16373 => x"30c30c",
   16374 => x"30c30c",
   16375 => x"30c30c",
   16376 => x"30c30c",
   16377 => x"30c30c",
   16378 => x"30c30c",
   16379 => x"30c30c",
   16380 => x"30c30c",
   16381 => x"30c30c",
   16382 => x"30c30c",
   16383 => x"30c30c",
   16384 => x"30c30c",
   16385 => x"30c30c",
   16386 => x"30c30c",
   16387 => x"30c30c",
   16388 => x"32efff",
   16389 => x"ffffff",
   16390 => x"ffffff",
   16391 => x"ffffff",
   16392 => x"ffffff",
   16393 => x"ffffff",
   16394 => x"ffffff",
   16395 => x"ffffff",
   16396 => x"ffffff",
   16397 => x"ffffff",
   16398 => x"ffffff",
   16399 => x"ffffff",
   16400 => x"ffffff",
   16401 => x"ffffff",
   16402 => x"ffffff",
   16403 => x"ffffff",
   16404 => x"ffffff",
   16405 => x"ffffff",
   16406 => x"a95abf",
   16407 => x"ffffff",
   16408 => x"ffffff",
   16409 => x"ffffff",
   16410 => x"ffffff",
   16411 => x"ffffff",
   16412 => x"ffffff",
   16413 => x"ffffff",
   16414 => x"ffffff",
   16415 => x"ffffff",
   16416 => x"ffffff",
   16417 => x"ffffff",
   16418 => x"ffffff",
   16419 => x"ffffff",
   16420 => x"ffffff",
   16421 => x"ffffff",
   16422 => x"ffffff",
   16423 => x"ffffff",
   16424 => x"ffffff",
   16425 => x"ffffff",
   16426 => x"ffffff",
   16427 => x"ffffff",
   16428 => x"ffffff",
   16429 => x"ffffff",
   16430 => x"ffffff",
   16431 => x"ffffff",
   16432 => x"ffffff",
   16433 => x"ffffff",
   16434 => x"ffffff",
   16435 => x"ffffff",
   16436 => x"ffffff",
   16437 => x"ffffff",
   16438 => x"ffffff",
   16439 => x"ffffff",
   16440 => x"ffffff",
   16441 => x"ffffff",
   16442 => x"ffffff",
   16443 => x"ffffff",
   16444 => x"ffffff",
   16445 => x"ffffff",
   16446 => x"ffffff",
   16447 => x"ffffff",
   16448 => x"ffffff",
   16449 => x"ffffff",
   16450 => x"ffffff",
   16451 => x"ffffff",
   16452 => x"ffffff",
   16453 => x"ffffff",
   16454 => x"ffffff",
   16455 => x"ffffff",
   16456 => x"ffffff",
   16457 => x"ffffff",
   16458 => x"ffffff",
   16459 => x"ffffff",
   16460 => x"ffffff",
   16461 => x"ffffff",
   16462 => x"ffffff",
   16463 => x"ffffff",
   16464 => x"ffffff",
   16465 => x"ffffff",
   16466 => x"ffffff",
   16467 => x"ffffff",
   16468 => x"ffffff",
   16469 => x"ffffff",
   16470 => x"ffffff",
   16471 => x"ffffff",
   16472 => x"ffffff",
   16473 => x"ffffff",
   16474 => x"ffffff",
   16475 => x"ffffff",
   16476 => x"ffffff",
   16477 => x"ffffff",
   16478 => x"ffffff",
   16479 => x"ffffff",
   16480 => x"ff5c30",
   16481 => x"c30c30",
   16482 => x"c30c30",
   16483 => x"c30c30",
   16484 => x"c30c30",
   16485 => x"c30c30",
   16486 => x"c30c30",
   16487 => x"c30c30",
   16488 => x"c30c30",
   16489 => x"c30c30",
   16490 => x"c30c30",
   16491 => x"c30c30",
   16492 => x"c30c30",
   16493 => x"c30c30",
   16494 => x"c30c30",
   16495 => x"c30c30",
   16496 => x"c30c30",
   16497 => x"c30c30",
   16498 => x"c30c30",
   16499 => x"c30c30",
   16500 => x"c30c30",
   16501 => x"c30c30",
   16502 => x"a2cf3c",
   16503 => x"f3cf3c",
   16504 => x"f3cf3c",
   16505 => x"f3cf3c",
   16506 => x"f3cf3c",
   16507 => x"f2cb1d",
   16508 => x"bbefff",
   16509 => x"ffffff",
   16510 => x"ffffff",
   16511 => x"ffffff",
   16512 => x"ffffff",
   16513 => x"ffffff",
   16514 => x"ffffff",
   16515 => x"ffffff",
   16516 => x"ffffff",
   16517 => x"ffffff",
   16518 => x"ffffff",
   16519 => x"ffffff",
   16520 => x"feeb9d",
   16521 => x"72cf3c",
   16522 => x"f3cf3c",
   16523 => x"f3cf3c",
   16524 => x"f3cf3c",
   16525 => x"f3cf3c",
   16526 => x"f2c30c",
   16527 => x"30c30c",
   16528 => x"30c30c",
   16529 => x"30c30c",
   16530 => x"30c30c",
   16531 => x"30c30c",
   16532 => x"30c30c",
   16533 => x"30c30c",
   16534 => x"30c30c",
   16535 => x"30c30c",
   16536 => x"30c30c",
   16537 => x"30c30c",
   16538 => x"30c30c",
   16539 => x"30c30c",
   16540 => x"30c30c",
   16541 => x"30c30c",
   16542 => x"30c30c",
   16543 => x"30c30c",
   16544 => x"30c30c",
   16545 => x"30c30c",
   16546 => x"30c30c",
   16547 => x"30c30c",
   16548 => x"32efff",
   16549 => x"ffffff",
   16550 => x"ffffff",
   16551 => x"ffffff",
   16552 => x"ffffff",
   16553 => x"ffffff",
   16554 => x"ffffff",
   16555 => x"ffffff",
   16556 => x"ffffff",
   16557 => x"ffffff",
   16558 => x"ffffff",
   16559 => x"ffffff",
   16560 => x"ffffff",
   16561 => x"ffffff",
   16562 => x"ffffff",
   16563 => x"ffffff",
   16564 => x"ffffff",
   16565 => x"ffffea",
   16566 => x"56afff",
   16567 => x"ffffff",
   16568 => x"ffffff",
   16569 => x"ffffff",
   16570 => x"ffffff",
   16571 => x"ffffff",
   16572 => x"ffffff",
   16573 => x"ffffff",
   16574 => x"ffffff",
   16575 => x"ffffff",
   16576 => x"ffffff",
   16577 => x"ffffff",
   16578 => x"ffffff",
   16579 => x"ffffff",
   16580 => x"ffffff",
   16581 => x"ffffff",
   16582 => x"ffffff",
   16583 => x"ffffff",
   16584 => x"ffffff",
   16585 => x"ffffff",
   16586 => x"ffffff",
   16587 => x"ffffff",
   16588 => x"ffffff",
   16589 => x"ffffff",
   16590 => x"ffffff",
   16591 => x"ffffff",
   16592 => x"ffffff",
   16593 => x"ffffff",
   16594 => x"ffffff",
   16595 => x"ffffff",
   16596 => x"ffffff",
   16597 => x"ffffff",
   16598 => x"ffffff",
   16599 => x"ffffff",
   16600 => x"ffffff",
   16601 => x"ffffff",
   16602 => x"ffffff",
   16603 => x"ffffff",
   16604 => x"ffffff",
   16605 => x"ffffff",
   16606 => x"ffffff",
   16607 => x"ffffff",
   16608 => x"ffffff",
   16609 => x"ffffff",
   16610 => x"ffffff",
   16611 => x"ffffff",
   16612 => x"ffffff",
   16613 => x"ffffff",
   16614 => x"ffffff",
   16615 => x"ffffff",
   16616 => x"ffffff",
   16617 => x"ffffff",
   16618 => x"ffffff",
   16619 => x"ffffff",
   16620 => x"ffffff",
   16621 => x"ffffff",
   16622 => x"ffffff",
   16623 => x"ffffff",
   16624 => x"ffffff",
   16625 => x"ffffff",
   16626 => x"ffffff",
   16627 => x"ffffff",
   16628 => x"ffffff",
   16629 => x"ffffff",
   16630 => x"ffffff",
   16631 => x"ffffff",
   16632 => x"ffffff",
   16633 => x"ffffff",
   16634 => x"ffffff",
   16635 => x"ffffff",
   16636 => x"ffffff",
   16637 => x"ffffff",
   16638 => x"ffffff",
   16639 => x"ffffff",
   16640 => x"ff5c30",
   16641 => x"c30c30",
   16642 => x"c30c30",
   16643 => x"c30c30",
   16644 => x"c30c30",
   16645 => x"c30c30",
   16646 => x"c30c30",
   16647 => x"c30c30",
   16648 => x"c30c30",
   16649 => x"c30c30",
   16650 => x"c30c30",
   16651 => x"c30c30",
   16652 => x"c30c30",
   16653 => x"c30c30",
   16654 => x"c30c30",
   16655 => x"c30c30",
   16656 => x"c30c30",
   16657 => x"c30c30",
   16658 => x"c30c30",
   16659 => x"c30c30",
   16660 => x"c30c30",
   16661 => x"c30c30",
   16662 => x"62cf3c",
   16663 => x"f3cf3c",
   16664 => x"f3cf3c",
   16665 => x"f3cf3c",
   16666 => x"f3cb1c",
   16667 => x"76efff",
   16668 => x"ffffff",
   16669 => x"ffffff",
   16670 => x"ffffff",
   16671 => x"ffffff",
   16672 => x"ffffff",
   16673 => x"ffffff",
   16674 => x"ffffff",
   16675 => x"ffffff",
   16676 => x"ffffff",
   16677 => x"ffffff",
   16678 => x"ffffff",
   16679 => x"ffffff",
   16680 => x"ffffff",
   16681 => x"fee75c",
   16682 => x"b3cf3c",
   16683 => x"f3cf3c",
   16684 => x"f3cf3c",
   16685 => x"f3cf3c",
   16686 => x"f2c30c",
   16687 => x"30c30c",
   16688 => x"30c30c",
   16689 => x"30c30c",
   16690 => x"30c30c",
   16691 => x"30c30c",
   16692 => x"30c30c",
   16693 => x"30c30c",
   16694 => x"30c30c",
   16695 => x"30c30c",
   16696 => x"30c30c",
   16697 => x"30c30c",
   16698 => x"30c30c",
   16699 => x"30c30c",
   16700 => x"30c30c",
   16701 => x"30c30c",
   16702 => x"30c30c",
   16703 => x"30c30c",
   16704 => x"30c30c",
   16705 => x"30c30c",
   16706 => x"30c30c",
   16707 => x"30c30c",
   16708 => x"32efff",
   16709 => x"ffffff",
   16710 => x"ffffff",
   16711 => x"ffffff",
   16712 => x"ffffff",
   16713 => x"ffffff",
   16714 => x"ffffff",
   16715 => x"ffffff",
   16716 => x"ffffff",
   16717 => x"ffffff",
   16718 => x"ffffff",
   16719 => x"ffffff",
   16720 => x"ffffff",
   16721 => x"ffffff",
   16722 => x"ffffff",
   16723 => x"ffffff",
   16724 => x"ffffff",
   16725 => x"fffa95",
   16726 => x"abffff",
   16727 => x"ffffff",
   16728 => x"ffffff",
   16729 => x"ffffff",
   16730 => x"ffffff",
   16731 => x"ffffff",
   16732 => x"ffffff",
   16733 => x"ffffff",
   16734 => x"ffffff",
   16735 => x"ffffff",
   16736 => x"ffffff",
   16737 => x"ffffff",
   16738 => x"ffffff",
   16739 => x"ffffff",
   16740 => x"ffffff",
   16741 => x"ffffff",
   16742 => x"ffffff",
   16743 => x"ffffff",
   16744 => x"ffffff",
   16745 => x"ffffff",
   16746 => x"ffffff",
   16747 => x"ffffff",
   16748 => x"ffffff",
   16749 => x"ffffff",
   16750 => x"ffffff",
   16751 => x"ffffff",
   16752 => x"ffffff",
   16753 => x"ffffff",
   16754 => x"ffffff",
   16755 => x"ffffff",
   16756 => x"ffffff",
   16757 => x"ffffff",
   16758 => x"ffffff",
   16759 => x"ffffff",
   16760 => x"ffffff",
   16761 => x"ffffff",
   16762 => x"ffffff",
   16763 => x"ffffff",
   16764 => x"ffffff",
   16765 => x"ffffff",
   16766 => x"ffffff",
   16767 => x"ffffff",
   16768 => x"ffffff",
   16769 => x"ffffff",
   16770 => x"ffffff",
   16771 => x"ffffff",
   16772 => x"ffffff",
   16773 => x"ffffff",
   16774 => x"ffffff",
   16775 => x"ffffff",
   16776 => x"ffffff",
   16777 => x"ffffff",
   16778 => x"ffffff",
   16779 => x"ffffff",
   16780 => x"ffffff",
   16781 => x"ffffff",
   16782 => x"ffffff",
   16783 => x"ffffff",
   16784 => x"ffffff",
   16785 => x"ffffff",
   16786 => x"ffffff",
   16787 => x"ffffff",
   16788 => x"ffffff",
   16789 => x"ffffff",
   16790 => x"ffffff",
   16791 => x"ffffff",
   16792 => x"ffffff",
   16793 => x"ffffff",
   16794 => x"ffffff",
   16795 => x"ffffff",
   16796 => x"ffffff",
   16797 => x"ffffff",
   16798 => x"ffffff",
   16799 => x"ffffff",
   16800 => x"ff5c30",
   16801 => x"c30c30",
   16802 => x"c30c30",
   16803 => x"c30c30",
   16804 => x"c30c30",
   16805 => x"c30c30",
   16806 => x"c30c30",
   16807 => x"c30c30",
   16808 => x"c30c30",
   16809 => x"c30c30",
   16810 => x"c30c30",
   16811 => x"c30c30",
   16812 => x"c30c30",
   16813 => x"c30c30",
   16814 => x"c30c30",
   16815 => x"c30c30",
   16816 => x"c30c30",
   16817 => x"c30c30",
   16818 => x"c30c30",
   16819 => x"c30c30",
   16820 => x"c30c30",
   16821 => x"c30c30",
   16822 => x"a2cf3c",
   16823 => x"f3cf3c",
   16824 => x"f3cf3c",
   16825 => x"f3cf2c",
   16826 => x"71dbbf",
   16827 => x"ffffff",
   16828 => x"ffffff",
   16829 => x"ffffff",
   16830 => x"ffffff",
   16831 => x"ffffff",
   16832 => x"ffffff",
   16833 => x"ffffff",
   16834 => x"ffffff",
   16835 => x"ffffff",
   16836 => x"ffffff",
   16837 => x"ffffff",
   16838 => x"ffffff",
   16839 => x"ffffff",
   16840 => x"ffffff",
   16841 => x"ffffff",
   16842 => x"b9d72c",
   16843 => x"f3cf3c",
   16844 => x"f3cf3c",
   16845 => x"f3cf3c",
   16846 => x"f2c30c",
   16847 => x"30c30c",
   16848 => x"30c30c",
   16849 => x"30c30c",
   16850 => x"30c30c",
   16851 => x"30c30c",
   16852 => x"30c30c",
   16853 => x"30c30c",
   16854 => x"30c30c",
   16855 => x"30c30c",
   16856 => x"30c30c",
   16857 => x"30c30c",
   16858 => x"30c30c",
   16859 => x"30c30c",
   16860 => x"30c30c",
   16861 => x"30c30c",
   16862 => x"30c30c",
   16863 => x"30c30c",
   16864 => x"30c30c",
   16865 => x"30c30c",
   16866 => x"30c30c",
   16867 => x"30c30c",
   16868 => x"32efff",
   16869 => x"ffffff",
   16870 => x"ffffff",
   16871 => x"ffffff",
   16872 => x"ffffff",
   16873 => x"ffffff",
   16874 => x"ffffff",
   16875 => x"ffffff",
   16876 => x"ffffff",
   16877 => x"ffffff",
   16878 => x"ffffff",
   16879 => x"ffffff",
   16880 => x"ffffff",
   16881 => x"ffffff",
   16882 => x"ffffff",
   16883 => x"ffffff",
   16884 => x"ffffff",
   16885 => x"fea56a",
   16886 => x"ffffff",
   16887 => x"ffffff",
   16888 => x"ffffff",
   16889 => x"ffffff",
   16890 => x"ffffff",
   16891 => x"ffffff",
   16892 => x"ffffff",
   16893 => x"ffffff",
   16894 => x"ffffff",
   16895 => x"ffffff",
   16896 => x"ffffff",
   16897 => x"ffffff",
   16898 => x"ffffff",
   16899 => x"ffffff",
   16900 => x"ffffff",
   16901 => x"ffffff",
   16902 => x"ffffff",
   16903 => x"ffffff",
   16904 => x"ffffff",
   16905 => x"ffffff",
   16906 => x"ffffff",
   16907 => x"ffffff",
   16908 => x"ffffff",
   16909 => x"ffffff",
   16910 => x"ffffff",
   16911 => x"ffffff",
   16912 => x"ffffff",
   16913 => x"ffffff",
   16914 => x"ffffff",
   16915 => x"ffffff",
   16916 => x"ffffff",
   16917 => x"ffffff",
   16918 => x"ffffff",
   16919 => x"ffffff",
   16920 => x"ffffff",
   16921 => x"ffffff",
   16922 => x"ffffff",
   16923 => x"ffffff",
   16924 => x"ffffff",
   16925 => x"ffffff",
   16926 => x"ffffff",
   16927 => x"ffffff",
   16928 => x"ffffff",
   16929 => x"ffffff",
   16930 => x"ffffff",
   16931 => x"ffffff",
   16932 => x"ffffff",
   16933 => x"ffffff",
   16934 => x"ffffff",
   16935 => x"ffffff",
   16936 => x"ffffff",
   16937 => x"ffffff",
   16938 => x"ffffff",
   16939 => x"ffffff",
   16940 => x"ffffff",
   16941 => x"ffffff",
   16942 => x"ffffff",
   16943 => x"ffffff",
   16944 => x"ffffff",
   16945 => x"ffffff",
   16946 => x"ffffff",
   16947 => x"ffffff",
   16948 => x"ffffff",
   16949 => x"ffffff",
   16950 => x"ffffff",
   16951 => x"ffffff",
   16952 => x"ffffff",
   16953 => x"ffffff",
   16954 => x"ffffff",
   16955 => x"ffffff",
   16956 => x"ffffff",
   16957 => x"ffffff",
   16958 => x"ffffff",
   16959 => x"ffffff",
   16960 => x"ff5c30",
   16961 => x"c30c30",
   16962 => x"c30c30",
   16963 => x"c30c30",
   16964 => x"c30c30",
   16965 => x"c30c30",
   16966 => x"c30c30",
   16967 => x"c30c30",
   16968 => x"c30c30",
   16969 => x"c30c30",
   16970 => x"c30c30",
   16971 => x"c30c30",
   16972 => x"c30c30",
   16973 => x"c30c30",
   16974 => x"c30c30",
   16975 => x"c30c30",
   16976 => x"c30c30",
   16977 => x"c30c30",
   16978 => x"c30c30",
   16979 => x"c30c30",
   16980 => x"c30c30",
   16981 => x"c30c30",
   16982 => x"a2cf3c",
   16983 => x"f3cf3c",
   16984 => x"f3cf3c",
   16985 => x"f2c71d",
   16986 => x"bbffff",
   16987 => x"ffffff",
   16988 => x"ffffff",
   16989 => x"ffffff",
   16990 => x"ffffff",
   16991 => x"ffffff",
   16992 => x"ffffff",
   16993 => x"ffffff",
   16994 => x"ffffff",
   16995 => x"ffffff",
   16996 => x"ffffff",
   16997 => x"ffffff",
   16998 => x"ffffff",
   16999 => x"ffffff",
   17000 => x"ffffff",
   17001 => x"ffffff",
   17002 => x"fffb9d",
   17003 => x"72cf3c",
   17004 => x"f3cf3c",
   17005 => x"f3cf3c",
   17006 => x"f2c30c",
   17007 => x"30c30c",
   17008 => x"30c30c",
   17009 => x"30c30c",
   17010 => x"30c30c",
   17011 => x"30c30c",
   17012 => x"30c30c",
   17013 => x"30c30c",
   17014 => x"30c30c",
   17015 => x"30c30c",
   17016 => x"30c30c",
   17017 => x"30c30c",
   17018 => x"30c30c",
   17019 => x"30c30c",
   17020 => x"30c30c",
   17021 => x"30c30c",
   17022 => x"30c30c",
   17023 => x"30c30c",
   17024 => x"30c30c",
   17025 => x"30c30c",
   17026 => x"30c30c",
   17027 => x"30c30c",
   17028 => x"32efff",
   17029 => x"ffffff",
   17030 => x"ffffff",
   17031 => x"ffffff",
   17032 => x"ffffff",
   17033 => x"ffffff",
   17034 => x"ffffff",
   17035 => x"ffffff",
   17036 => x"ffffff",
   17037 => x"ffffff",
   17038 => x"ffffff",
   17039 => x"ffffff",
   17040 => x"ffffff",
   17041 => x"ffffff",
   17042 => x"ffffff",
   17043 => x"ffffff",
   17044 => x"ffffff",
   17045 => x"a95abf",
   17046 => x"ffffff",
   17047 => x"ffffff",
   17048 => x"ffffff",
   17049 => x"ffffff",
   17050 => x"ffffff",
   17051 => x"ffffff",
   17052 => x"ffffff",
   17053 => x"ffffff",
   17054 => x"ffffff",
   17055 => x"ffffff",
   17056 => x"ffffff",
   17057 => x"ffffff",
   17058 => x"ffffff",
   17059 => x"ffffff",
   17060 => x"ffffff",
   17061 => x"ffffff",
   17062 => x"ffffff",
   17063 => x"ffffff",
   17064 => x"ffffff",
   17065 => x"ffffff",
   17066 => x"ffffff",
   17067 => x"ffffff",
   17068 => x"ffffff",
   17069 => x"ffffff",
   17070 => x"ffffff",
   17071 => x"ffffff",
   17072 => x"ffffff",
   17073 => x"ffffff",
   17074 => x"ffffff",
   17075 => x"ffffff",
   17076 => x"ffffff",
   17077 => x"ffffff",
   17078 => x"ffffff",
   17079 => x"ffffff",
   17080 => x"ffffff",
   17081 => x"ffffff",
   17082 => x"ffffff",
   17083 => x"ffffff",
   17084 => x"ffffff",
   17085 => x"ffffff",
   17086 => x"ffffff",
   17087 => x"ffffff",
   17088 => x"ffffff",
   17089 => x"ffffff",
   17090 => x"ffffff",
   17091 => x"ffffff",
   17092 => x"ffffff",
   17093 => x"ffffff",
   17094 => x"ffffff",
   17095 => x"ffffff",
   17096 => x"ffffff",
   17097 => x"ffffff",
   17098 => x"ffffff",
   17099 => x"ffffff",
   17100 => x"ffffff",
   17101 => x"ffffff",
   17102 => x"ffffff",
   17103 => x"ffffff",
   17104 => x"ffffff",
   17105 => x"ffffff",
   17106 => x"ffffff",
   17107 => x"ffffff",
   17108 => x"ffffff",
   17109 => x"ffffff",
   17110 => x"ffffff",
   17111 => x"ffffff",
   17112 => x"ffffff",
   17113 => x"ffffff",
   17114 => x"ffffff",
   17115 => x"ffffff",
   17116 => x"ffffff",
   17117 => x"ffffff",
   17118 => x"ffffff",
   17119 => x"ffffff",
   17120 => x"ff5c30",
   17121 => x"c30c30",
   17122 => x"c30c30",
   17123 => x"c30c30",
   17124 => x"c30c30",
   17125 => x"c30c30",
   17126 => x"c30c30",
   17127 => x"c30c30",
   17128 => x"c30c30",
   17129 => x"c30c30",
   17130 => x"c30c30",
   17131 => x"c30c30",
   17132 => x"c30c30",
   17133 => x"c30c30",
   17134 => x"c30c30",
   17135 => x"c30c30",
   17136 => x"c30c30",
   17137 => x"c30c30",
   17138 => x"c30c30",
   17139 => x"c30c30",
   17140 => x"c30c30",
   17141 => x"c30c30",
   17142 => x"92cf3c",
   17143 => x"f3cf3c",
   17144 => x"f3cb1c",
   17145 => x"76efff",
   17146 => x"ffffff",
   17147 => x"ffffff",
   17148 => x"ffffff",
   17149 => x"ffffff",
   17150 => x"ffffff",
   17151 => x"ffffff",
   17152 => x"ffffff",
   17153 => x"ffffff",
   17154 => x"ffffff",
   17155 => x"ffffff",
   17156 => x"ffffff",
   17157 => x"ffffff",
   17158 => x"ffffff",
   17159 => x"ffffff",
   17160 => x"ffffff",
   17161 => x"ffffff",
   17162 => x"ffffff",
   17163 => x"bae75c",
   17164 => x"b3cf3c",
   17165 => x"f3cf3c",
   17166 => x"f2c30c",
   17167 => x"30c30c",
   17168 => x"30c30c",
   17169 => x"30c30c",
   17170 => x"30c30c",
   17171 => x"30c30c",
   17172 => x"30c30c",
   17173 => x"30c30c",
   17174 => x"30c30c",
   17175 => x"30c30c",
   17176 => x"30c30c",
   17177 => x"30c30c",
   17178 => x"30c30c",
   17179 => x"30c30c",
   17180 => x"30c30c",
   17181 => x"30c30c",
   17182 => x"30c30c",
   17183 => x"30c30c",
   17184 => x"30c30c",
   17185 => x"30c30c",
   17186 => x"30c30c",
   17187 => x"30c30c",
   17188 => x"32efff",
   17189 => x"ffffff",
   17190 => x"ffffff",
   17191 => x"ffffff",
   17192 => x"ffffff",
   17193 => x"ffffff",
   17194 => x"ffffff",
   17195 => x"ffffff",
   17196 => x"ffffff",
   17197 => x"ffffff",
   17198 => x"ffffff",
   17199 => x"ffffff",
   17200 => x"ffffff",
   17201 => x"ffffff",
   17202 => x"ffffff",
   17203 => x"ffffff",
   17204 => x"ffffea",
   17205 => x"56afff",
   17206 => x"ffffff",
   17207 => x"ffffff",
   17208 => x"ffffff",
   17209 => x"ffffff",
   17210 => x"ffffff",
   17211 => x"ffffff",
   17212 => x"ffffff",
   17213 => x"ffffff",
   17214 => x"ffffff",
   17215 => x"ffffff",
   17216 => x"ffffff",
   17217 => x"ffffff",
   17218 => x"ffffff",
   17219 => x"ffffff",
   17220 => x"ffffff",
   17221 => x"ffffff",
   17222 => x"ffffff",
   17223 => x"ffffff",
   17224 => x"ffffff",
   17225 => x"ffffff",
   17226 => x"ffffff",
   17227 => x"ffffff",
   17228 => x"ffffff",
   17229 => x"ffffff",
   17230 => x"ffffff",
   17231 => x"ffffff",
   17232 => x"ffffff",
   17233 => x"ffffff",
   17234 => x"ffffff",
   17235 => x"ffffff",
   17236 => x"ffffff",
   17237 => x"ffffff",
   17238 => x"ffffff",
   17239 => x"ffffff",
   17240 => x"ffffff",
   17241 => x"ffffff",
   17242 => x"ffffff",
   17243 => x"ffffff",
   17244 => x"ffffff",
   17245 => x"ffffff",
   17246 => x"ffffff",
   17247 => x"ffffff",
   17248 => x"ffffff",
   17249 => x"ffffff",
   17250 => x"ffffff",
   17251 => x"ffffff",
   17252 => x"ffffff",
   17253 => x"ffffff",
   17254 => x"ffffff",
   17255 => x"ffffff",
   17256 => x"ffffff",
   17257 => x"ffffff",
   17258 => x"ffffff",
   17259 => x"ffffff",
   17260 => x"ffffff",
   17261 => x"ffffff",
   17262 => x"ffffff",
   17263 => x"ffffff",
   17264 => x"ffffff",
   17265 => x"ffffff",
   17266 => x"ffffff",
   17267 => x"ffffff",
   17268 => x"ffffff",
   17269 => x"ffffff",
   17270 => x"ffffff",
   17271 => x"ffffff",
   17272 => x"ffffff",
   17273 => x"ffffff",
   17274 => x"ffffff",
   17275 => x"ffffff",
   17276 => x"ffffff",
   17277 => x"ffffff",
   17278 => x"ffffff",
   17279 => x"ffffff",
   17280 => x"ff5c30",
   17281 => x"c30c30",
   17282 => x"c30c30",
   17283 => x"c30c30",
   17284 => x"c30c30",
   17285 => x"c30c30",
   17286 => x"c30c30",
   17287 => x"c30c30",
   17288 => x"c30c30",
   17289 => x"c30c30",
   17290 => x"c30c30",
   17291 => x"c30c30",
   17292 => x"c30c30",
   17293 => x"c30c30",
   17294 => x"c30c30",
   17295 => x"c30c30",
   17296 => x"c30c30",
   17297 => x"c30c30",
   17298 => x"c30c30",
   17299 => x"c30c30",
   17300 => x"c30c30",
   17301 => x"c30c30",
   17302 => x"92cf3c",
   17303 => x"f3cf3c",
   17304 => x"b1c76e",
   17305 => x"ffffff",
   17306 => x"ffffff",
   17307 => x"ffffff",
   17308 => x"ffffff",
   17309 => x"ffffff",
   17310 => x"ffffff",
   17311 => x"ffffff",
   17312 => x"ffffff",
   17313 => x"ffffff",
   17314 => x"ffffff",
   17315 => x"ffffff",
   17316 => x"ffffff",
   17317 => x"ffffff",
   17318 => x"ffffff",
   17319 => x"ffffff",
   17320 => x"ffffff",
   17321 => x"ffffff",
   17322 => x"ffffff",
   17323 => x"ffffee",
   17324 => x"75cb3c",
   17325 => x"f3cf3c",
   17326 => x"f2c30c",
   17327 => x"30c30c",
   17328 => x"30c30c",
   17329 => x"30c30c",
   17330 => x"30c30c",
   17331 => x"30c30c",
   17332 => x"30c30c",
   17333 => x"30c30c",
   17334 => x"30c30c",
   17335 => x"30c30c",
   17336 => x"30c30c",
   17337 => x"30c30c",
   17338 => x"30c30c",
   17339 => x"30c30c",
   17340 => x"30c30c",
   17341 => x"30c30c",
   17342 => x"30c30c",
   17343 => x"30c30c",
   17344 => x"30c30c",
   17345 => x"30c30c",
   17346 => x"30c30c",
   17347 => x"30c30c",
   17348 => x"32efff",
   17349 => x"ffffff",
   17350 => x"ffffff",
   17351 => x"ffffff",
   17352 => x"ffffff",
   17353 => x"ffffff",
   17354 => x"ffffff",
   17355 => x"ffffff",
   17356 => x"ffffff",
   17357 => x"ffffff",
   17358 => x"ffffff",
   17359 => x"ffffff",
   17360 => x"ffffff",
   17361 => x"ffffff",
   17362 => x"ffffff",
   17363 => x"ffffff",
   17364 => x"fffa95",
   17365 => x"abffff",
   17366 => x"ffffff",
   17367 => x"ffffff",
   17368 => x"ffffff",
   17369 => x"ffffff",
   17370 => x"ffffff",
   17371 => x"ffffff",
   17372 => x"ffffff",
   17373 => x"ffffff",
   17374 => x"ffffff",
   17375 => x"ffffff",
   17376 => x"ffffff",
   17377 => x"ffffff",
   17378 => x"ffffff",
   17379 => x"ffffff",
   17380 => x"ffffff",
   17381 => x"ffffff",
   17382 => x"ffffff",
   17383 => x"ffffff",
   17384 => x"ffffff",
   17385 => x"ffffff",
   17386 => x"ffffff",
   17387 => x"ffffff",
   17388 => x"ffffff",
   17389 => x"ffffff",
   17390 => x"ffffff",
   17391 => x"ffffff",
   17392 => x"ffffff",
   17393 => x"ffffff",
   17394 => x"ffffff",
   17395 => x"ffffff",
   17396 => x"ffffff",
   17397 => x"ffffff",
   17398 => x"ffffff",
   17399 => x"ffffff",
   17400 => x"ffffff",
   17401 => x"ffffff",
   17402 => x"ffffff",
   17403 => x"ffffff",
   17404 => x"ffffff",
   17405 => x"ffffff",
   17406 => x"ffffff",
   17407 => x"ffffff",
   17408 => x"ffffff",
   17409 => x"ffffff",
   17410 => x"ffffff",
   17411 => x"ffffff",
   17412 => x"ffffff",
   17413 => x"ffffff",
   17414 => x"ffffff",
   17415 => x"ffffff",
   17416 => x"ffffff",
   17417 => x"ffffff",
   17418 => x"ffffff",
   17419 => x"ffffff",
   17420 => x"ffffff",
   17421 => x"ffffff",
   17422 => x"ffffff",
   17423 => x"ffffff",
   17424 => x"ffffff",
   17425 => x"ffffff",
   17426 => x"ffffff",
   17427 => x"ffffff",
   17428 => x"ffffff",
   17429 => x"ffffff",
   17430 => x"ffffff",
   17431 => x"ffffff",
   17432 => x"ffffff",
   17433 => x"ffffff",
   17434 => x"ffffff",
   17435 => x"ffffff",
   17436 => x"ffffff",
   17437 => x"ffffff",
   17438 => x"ffffff",
   17439 => x"ffffff",
   17440 => x"ff5c30",
   17441 => x"c30c30",
   17442 => x"c30c30",
   17443 => x"c30c30",
   17444 => x"c30c30",
   17445 => x"c30c30",
   17446 => x"c30c30",
   17447 => x"c30c30",
   17448 => x"c30c30",
   17449 => x"c30c30",
   17450 => x"c30c30",
   17451 => x"c30c30",
   17452 => x"c30c30",
   17453 => x"c30c30",
   17454 => x"c30c30",
   17455 => x"c30c30",
   17456 => x"c30c30",
   17457 => x"c30c30",
   17458 => x"c30c30",
   17459 => x"c30c30",
   17460 => x"c30c30",
   17461 => x"c30c30",
   17462 => x"92cf3c",
   17463 => x"f3cb1d",
   17464 => x"bbefff",
   17465 => x"ffffff",
   17466 => x"ffffff",
   17467 => x"ffffff",
   17468 => x"ffffff",
   17469 => x"ffffff",
   17470 => x"ffffff",
   17471 => x"ffffff",
   17472 => x"ffffff",
   17473 => x"ffffff",
   17474 => x"ffffff",
   17475 => x"ffffff",
   17476 => x"ffffff",
   17477 => x"ffffff",
   17478 => x"ffffff",
   17479 => x"ffffff",
   17480 => x"ffffff",
   17481 => x"ffffff",
   17482 => x"ffffff",
   17483 => x"ffffff",
   17484 => x"feeb5c",
   17485 => x"b3cf3c",
   17486 => x"f2c30c",
   17487 => x"30c30c",
   17488 => x"30c30c",
   17489 => x"30c30c",
   17490 => x"30c30c",
   17491 => x"30c30c",
   17492 => x"30c30c",
   17493 => x"30c30c",
   17494 => x"30c30c",
   17495 => x"30c30c",
   17496 => x"30c30c",
   17497 => x"30c30c",
   17498 => x"30c30c",
   17499 => x"30c30c",
   17500 => x"30c30c",
   17501 => x"30c30c",
   17502 => x"30c30c",
   17503 => x"30c30c",
   17504 => x"30c30c",
   17505 => x"30c30c",
   17506 => x"30c30c",
   17507 => x"30c30c",
   17508 => x"32efff",
   17509 => x"ffffff",
   17510 => x"ffffff",
   17511 => x"ffffff",
   17512 => x"ffffff",
   17513 => x"ffffff",
   17514 => x"ffffff",
   17515 => x"ffffff",
   17516 => x"ffffff",
   17517 => x"ffffff",
   17518 => x"ffffff",
   17519 => x"ffffff",
   17520 => x"ffffff",
   17521 => x"ffffff",
   17522 => x"ffffff",
   17523 => x"ffffff",
   17524 => x"fea56a",
   17525 => x"ffffff",
   17526 => x"ffffff",
   17527 => x"ffffff",
   17528 => x"ffffff",
   17529 => x"ffffff",
   17530 => x"ffffff",
   17531 => x"ffffff",
   17532 => x"ffffff",
   17533 => x"ffffff",
   17534 => x"ffffff",
   17535 => x"ffffff",
   17536 => x"ffffff",
   17537 => x"ffffff",
   17538 => x"ffffff",
   17539 => x"ffffff",
   17540 => x"ffffff",
   17541 => x"ffffff",
   17542 => x"ffffff",
   17543 => x"ffffff",
   17544 => x"ffffff",
   17545 => x"ffffff",
   17546 => x"ffffff",
   17547 => x"ffffff",
   17548 => x"ffffff",
   17549 => x"ffffff",
   17550 => x"ffffff",
   17551 => x"ffffff",
   17552 => x"ffffff",
   17553 => x"ffffff",
   17554 => x"ffffff",
   17555 => x"ffffff",
   17556 => x"ffffff",
   17557 => x"ffffff",
   17558 => x"ffffff",
   17559 => x"ffffff",
   17560 => x"ffffff",
   17561 => x"ffffff",
   17562 => x"ffffff",
   17563 => x"ffffff",
   17564 => x"ffffff",
   17565 => x"ffffff",
   17566 => x"ffffff",
   17567 => x"ffffff",
   17568 => x"ffffff",
   17569 => x"ffffff",
   17570 => x"ffffff",
   17571 => x"ffffff",
   17572 => x"ffffff",
   17573 => x"ffffff",
   17574 => x"ffffff",
   17575 => x"ffffff",
   17576 => x"ffffff",
   17577 => x"ffffff",
   17578 => x"ffffff",
   17579 => x"ffffff",
   17580 => x"ffffff",
   17581 => x"ffffff",
   17582 => x"ffffff",
   17583 => x"ffffff",
   17584 => x"ffffff",
   17585 => x"ffffff",
   17586 => x"ffffff",
   17587 => x"ffffff",
   17588 => x"ffffff",
   17589 => x"ffffff",
   17590 => x"ffffff",
   17591 => x"ffffff",
   17592 => x"ffffff",
   17593 => x"ffffff",
   17594 => x"ffffff",
   17595 => x"ffffff",
   17596 => x"ffffff",
   17597 => x"ffffff",
   17598 => x"ffffff",
   17599 => x"ffffff",
   17600 => x"ffac30",
   17601 => x"c30c30",
   17602 => x"c30c30",
   17603 => x"c30c30",
   17604 => x"c30c30",
   17605 => x"c30c30",
   17606 => x"c30c30",
   17607 => x"c30c30",
   17608 => x"c30c30",
   17609 => x"c30c30",
   17610 => x"c30c30",
   17611 => x"c30c30",
   17612 => x"c30c30",
   17613 => x"c30c30",
   17614 => x"c30c30",
   17615 => x"c30c30",
   17616 => x"c30c30",
   17617 => x"c30c30",
   17618 => x"c30c30",
   17619 => x"c30c30",
   17620 => x"c30c30",
   17621 => x"c30c30",
   17622 => x"92cf3c",
   17623 => x"b1cbae",
   17624 => x"ffffff",
   17625 => x"ffffff",
   17626 => x"ffffff",
   17627 => x"ffffff",
   17628 => x"ffffff",
   17629 => x"ffffff",
   17630 => x"ffffff",
   17631 => x"ffffff",
   17632 => x"ffffff",
   17633 => x"ffffff",
   17634 => x"ffffff",
   17635 => x"ffffff",
   17636 => x"ffffff",
   17637 => x"ffffff",
   17638 => x"ffffff",
   17639 => x"ffffff",
   17640 => x"ffffff",
   17641 => x"ffffff",
   17642 => x"ffffff",
   17643 => x"ffffff",
   17644 => x"ffffee",
   17645 => x"b5cb3c",
   17646 => x"f2c30c",
   17647 => x"30c30c",
   17648 => x"30c30c",
   17649 => x"30c30c",
   17650 => x"30c30c",
   17651 => x"30c30c",
   17652 => x"30c30c",
   17653 => x"30c30c",
   17654 => x"30c30c",
   17655 => x"30c30c",
   17656 => x"30c30c",
   17657 => x"30c30c",
   17658 => x"30c30c",
   17659 => x"30c30c",
   17660 => x"30c30c",
   17661 => x"30c30c",
   17662 => x"30c30c",
   17663 => x"30c30c",
   17664 => x"30c30c",
   17665 => x"30c30c",
   17666 => x"30c30c",
   17667 => x"30c30c",
   17668 => x"32efff",
   17669 => x"ffffff",
   17670 => x"ffffff",
   17671 => x"ffffff",
   17672 => x"ffffff",
   17673 => x"ffffff",
   17674 => x"ffffff",
   17675 => x"ffffff",
   17676 => x"ffffff",
   17677 => x"ffffff",
   17678 => x"ffffff",
   17679 => x"ffffff",
   17680 => x"ffffff",
   17681 => x"ffffff",
   17682 => x"ffffff",
   17683 => x"ffffff",
   17684 => x"a95abf",
   17685 => x"ffffff",
   17686 => x"ffffff",
   17687 => x"ffffff",
   17688 => x"ffffff",
   17689 => x"ffffff",
   17690 => x"ffffff",
   17691 => x"ffffff",
   17692 => x"ffffff",
   17693 => x"ffffff",
   17694 => x"ffffff",
   17695 => x"ffffff",
   17696 => x"ffffff",
   17697 => x"ffffff",
   17698 => x"ffffff",
   17699 => x"ffffff",
   17700 => x"ffffff",
   17701 => x"ffffff",
   17702 => x"ffffff",
   17703 => x"ffffff",
   17704 => x"ffffff",
   17705 => x"ffffff",
   17706 => x"ffffff",
   17707 => x"ffffff",
   17708 => x"ffffff",
   17709 => x"ffffff",
   17710 => x"ffffff",
   17711 => x"ffffff",
   17712 => x"ffffff",
   17713 => x"ffffff",
   17714 => x"ffffff",
   17715 => x"ffffff",
   17716 => x"ffffff",
   17717 => x"ffffff",
   17718 => x"ffffff",
   17719 => x"ffffff",
   17720 => x"ffffff",
   17721 => x"ffffff",
   17722 => x"ffffff",
   17723 => x"ffffff",
   17724 => x"ffffff",
   17725 => x"ffffff",
   17726 => x"ffffff",
   17727 => x"ffffff",
   17728 => x"ffffff",
   17729 => x"ffffff",
   17730 => x"ffffff",
   17731 => x"ffffff",
   17732 => x"ffffff",
   17733 => x"ffffff",
   17734 => x"ffffff",
   17735 => x"ffffff",
   17736 => x"ffffff",
   17737 => x"ffffff",
   17738 => x"ffffff",
   17739 => x"ffffff",
   17740 => x"ffffff",
   17741 => x"ffffff",
   17742 => x"ffffff",
   17743 => x"ffffff",
   17744 => x"ffffff",
   17745 => x"ffffff",
   17746 => x"ffffff",
   17747 => x"ffffff",
   17748 => x"ffffff",
   17749 => x"ffffff",
   17750 => x"ffffff",
   17751 => x"ffffff",
   17752 => x"ffffff",
   17753 => x"ffffff",
   17754 => x"ffffff",
   17755 => x"ffffff",
   17756 => x"ffffff",
   17757 => x"ffffff",
   17758 => x"ffffff",
   17759 => x"ffffff",
   17760 => x"ffac30",
   17761 => x"c30c30",
   17762 => x"c30c30",
   17763 => x"c30c30",
   17764 => x"c30c30",
   17765 => x"c30c30",
   17766 => x"c30c30",
   17767 => x"c30c30",
   17768 => x"c30c30",
   17769 => x"c30c30",
   17770 => x"c30c30",
   17771 => x"c30c30",
   17772 => x"c30c30",
   17773 => x"c30c30",
   17774 => x"c30c30",
   17775 => x"c30c30",
   17776 => x"c30c30",
   17777 => x"c30c30",
   17778 => x"c30c30",
   17779 => x"c30c30",
   17780 => x"c30c30",
   17781 => x"c30c30",
   17782 => x"92cb1c",
   17783 => x"b6efff",
   17784 => x"ffffff",
   17785 => x"ffffff",
   17786 => x"ffffff",
   17787 => x"ffffff",
   17788 => x"ffffff",
   17789 => x"ffffff",
   17790 => x"ffffff",
   17791 => x"ffffff",
   17792 => x"ffffff",
   17793 => x"ffffff",
   17794 => x"ffffff",
   17795 => x"ffffff",
   17796 => x"ffffff",
   17797 => x"ffffff",
   17798 => x"ffffff",
   17799 => x"ffffff",
   17800 => x"ffffff",
   17801 => x"ffffff",
   17802 => x"ffffff",
   17803 => x"ffffff",
   17804 => x"ffffff",
   17805 => x"fee75c",
   17806 => x"b2c30c",
   17807 => x"30c30c",
   17808 => x"30c30c",
   17809 => x"30c30c",
   17810 => x"30c30c",
   17811 => x"30c30c",
   17812 => x"30c30c",
   17813 => x"30c30c",
   17814 => x"30c30c",
   17815 => x"30c30c",
   17816 => x"30c30c",
   17817 => x"30c30c",
   17818 => x"30c30c",
   17819 => x"30c30c",
   17820 => x"30c30c",
   17821 => x"30c30c",
   17822 => x"30c30c",
   17823 => x"30c30c",
   17824 => x"30c30c",
   17825 => x"30c30c",
   17826 => x"30c30c",
   17827 => x"30c30c",
   17828 => x"76efff",
   17829 => x"ffffff",
   17830 => x"ffffff",
   17831 => x"ffffff",
   17832 => x"ffffff",
   17833 => x"ffffff",
   17834 => x"ffffff",
   17835 => x"ffffff",
   17836 => x"ffffff",
   17837 => x"ffffff",
   17838 => x"ffffff",
   17839 => x"ffffff",
   17840 => x"ffffff",
   17841 => x"ffffff",
   17842 => x"ffffff",
   17843 => x"ffffea",
   17844 => x"56afff",
   17845 => x"ffffff",
   17846 => x"ffffff",
   17847 => x"ffffff",
   17848 => x"ffffff",
   17849 => x"ffffff",
   17850 => x"ffffff",
   17851 => x"ffffff",
   17852 => x"ffffff",
   17853 => x"ffffff",
   17854 => x"ffffff",
   17855 => x"ffffff",
   17856 => x"ffffff",
   17857 => x"ffffff",
   17858 => x"ffffff",
   17859 => x"ffffff",
   17860 => x"ffffff",
   17861 => x"ffffff",
   17862 => x"ffffff",
   17863 => x"ffffff",
   17864 => x"ffffff",
   17865 => x"ffffff",
   17866 => x"ffffff",
   17867 => x"ffffff",
   17868 => x"ffffff",
   17869 => x"ffffff",
   17870 => x"ffffff",
   17871 => x"ffffff",
   17872 => x"ffffff",
   17873 => x"ffffff",
   17874 => x"ffffff",
   17875 => x"ffffff",
   17876 => x"ffffff",
   17877 => x"ffffff",
   17878 => x"ffffff",
   17879 => x"ffffff",
   17880 => x"ffffff",
   17881 => x"ffffff",
   17882 => x"ffffff",
   17883 => x"ffffff",
   17884 => x"ffffff",
   17885 => x"ffffff",
   17886 => x"ffffff",
   17887 => x"ffffff",
   17888 => x"ffffff",
   17889 => x"ffffff",
   17890 => x"ffffff",
   17891 => x"ffffff",
   17892 => x"ffffff",
   17893 => x"ffffff",
   17894 => x"ffffff",
   17895 => x"ffffff",
   17896 => x"ffffff",
   17897 => x"ffffff",
   17898 => x"ffffff",
   17899 => x"ffffff",
   17900 => x"ffffff",
   17901 => x"ffffff",
   17902 => x"ffffff",
   17903 => x"ffffff",
   17904 => x"ffffff",
   17905 => x"ffffff",
   17906 => x"ffffff",
   17907 => x"ffffff",
   17908 => x"ffffff",
   17909 => x"ffffff",
   17910 => x"ffffff",
   17911 => x"ffffff",
   17912 => x"ffffff",
   17913 => x"ffffff",
   17914 => x"ffffff",
   17915 => x"ffffff",
   17916 => x"ffffff",
   17917 => x"ffffff",
   17918 => x"ffffff",
   17919 => x"ffffff",
   17920 => x"ffac30",
   17921 => x"c30c30",
   17922 => x"c30c30",
   17923 => x"c30c30",
   17924 => x"c30c30",
   17925 => x"c30c30",
   17926 => x"c30c30",
   17927 => x"c30c30",
   17928 => x"c30c30",
   17929 => x"c30c30",
   17930 => x"c30c30",
   17931 => x"c30c30",
   17932 => x"c30c30",
   17933 => x"c30c30",
   17934 => x"c30c30",
   17935 => x"c30c30",
   17936 => x"c30c30",
   17937 => x"c30c30",
   17938 => x"c30c30",
   17939 => x"c30c30",
   17940 => x"c30c30",
   17941 => x"c30c30",
   17942 => x"91876e",
   17943 => x"ffffff",
   17944 => x"ffffff",
   17945 => x"ffffff",
   17946 => x"ffffff",
   17947 => x"ffffff",
   17948 => x"ffffff",
   17949 => x"ffffff",
   17950 => x"ffffff",
   17951 => x"ffffff",
   17952 => x"ffffff",
   17953 => x"ffffff",
   17954 => x"ffffff",
   17955 => x"ffffff",
   17956 => x"ffffff",
   17957 => x"ffffff",
   17958 => x"ffffff",
   17959 => x"ffffff",
   17960 => x"ffffff",
   17961 => x"ffffff",
   17962 => x"ffffff",
   17963 => x"ffffff",
   17964 => x"ffffff",
   17965 => x"ffffee",
   17966 => x"70c30c",
   17967 => x"30c30c",
   17968 => x"30c30c",
   17969 => x"30c30c",
   17970 => x"30c30c",
   17971 => x"30c30c",
   17972 => x"30c30c",
   17973 => x"30c30c",
   17974 => x"30c30c",
   17975 => x"30c30c",
   17976 => x"30c30c",
   17977 => x"30c30c",
   17978 => x"30c30c",
   17979 => x"30c30c",
   17980 => x"30c30c",
   17981 => x"30c30c",
   17982 => x"30c30c",
   17983 => x"30c30c",
   17984 => x"30c30c",
   17985 => x"30c30c",
   17986 => x"30c30c",
   17987 => x"30c30c",
   17988 => x"76efff",
   17989 => x"ffffff",
   17990 => x"ffffff",
   17991 => x"ffffff",
   17992 => x"ffffff",
   17993 => x"ffffff",
   17994 => x"ffffff",
   17995 => x"ffffff",
   17996 => x"ffffff",
   17997 => x"ffffff",
   17998 => x"ffffff",
   17999 => x"ffffff",
   18000 => x"ffffff",
   18001 => x"ffffff",
   18002 => x"ffffff",
   18003 => x"fffa95",
   18004 => x"abffff",
   18005 => x"ffffff",
   18006 => x"ffffff",
   18007 => x"ffffff",
   18008 => x"ffffff",
   18009 => x"ffffff",
   18010 => x"ffffff",
   18011 => x"ffffff",
   18012 => x"ffffff",
   18013 => x"ffffff",
   18014 => x"ffffff",
   18015 => x"ffffff",
   18016 => x"ffffff",
   18017 => x"ffffff",
   18018 => x"ffffff",
   18019 => x"ffffff",
   18020 => x"ffffff",
   18021 => x"ffffff",
   18022 => x"ffffff",
   18023 => x"ffffff",
   18024 => x"ffffff",
   18025 => x"ffffff",
   18026 => x"ffffff",
   18027 => x"ffffff",
   18028 => x"ffffff",
   18029 => x"ffffff",
   18030 => x"ffffff",
   18031 => x"ffffff",
   18032 => x"ffffff",
   18033 => x"ffffff",
   18034 => x"ffffff",
   18035 => x"ffffff",
   18036 => x"ffffff",
   18037 => x"ffffff",
   18038 => x"ffffff",
   18039 => x"ffffff",
   18040 => x"ffffff",
   18041 => x"ffffff",
   18042 => x"ffffff",
   18043 => x"ffffff",
   18044 => x"ffffff",
   18045 => x"ffffff",
   18046 => x"ffffff",
   18047 => x"ffffff",
   18048 => x"ffffff",
   18049 => x"ffffff",
   18050 => x"ffffff",
   18051 => x"ffffff",
   18052 => x"ffffff",
   18053 => x"ffffff",
   18054 => x"ffffff",
   18055 => x"ffffff",
   18056 => x"ffffff",
   18057 => x"ffffff",
   18058 => x"ffffff",
   18059 => x"ffffff",
   18060 => x"ffffff",
   18061 => x"ffffff",
   18062 => x"ffffff",
   18063 => x"ffffff",
   18064 => x"ffffff",
   18065 => x"ffffff",
   18066 => x"ffffff",
   18067 => x"ffffff",
   18068 => x"ffffff",
   18069 => x"ffffff",
   18070 => x"ffffff",
   18071 => x"ffffff",
   18072 => x"ffffff",
   18073 => x"ffffff",
   18074 => x"ffffff",
   18075 => x"ffffff",
   18076 => x"ffffff",
   18077 => x"ffffff",
   18078 => x"ffffff",
   18079 => x"ffffff",
   18080 => x"ffac30",
   18081 => x"c30c30",
   18082 => x"c30c30",
   18083 => x"c30c30",
   18084 => x"c30c30",
   18085 => x"c30c30",
   18086 => x"c30c30",
   18087 => x"c30c30",
   18088 => x"c30c30",
   18089 => x"c30c30",
   18090 => x"c30c30",
   18091 => x"c30c30",
   18092 => x"c30c30",
   18093 => x"c30c30",
   18094 => x"c30c30",
   18095 => x"c30c30",
   18096 => x"c30c30",
   18097 => x"c30c30",
   18098 => x"c30c30",
   18099 => x"c30c30",
   18100 => x"c30c30",
   18101 => x"c30c21",
   18102 => x"55abbf",
   18103 => x"ffffff",
   18104 => x"ffffff",
   18105 => x"ffffff",
   18106 => x"ffffff",
   18107 => x"ffffff",
   18108 => x"ffffff",
   18109 => x"ffffff",
   18110 => x"ffffff",
   18111 => x"ffffff",
   18112 => x"ffffff",
   18113 => x"ffffff",
   18114 => x"ffffff",
   18115 => x"ffffff",
   18116 => x"ffffff",
   18117 => x"ffffff",
   18118 => x"ffffff",
   18119 => x"ffffff",
   18120 => x"ffffff",
   18121 => x"ffffff",
   18122 => x"ffffff",
   18123 => x"ffffff",
   18124 => x"ffffff",
   18125 => x"ffffff",
   18126 => x"b8c34c",
   18127 => x"30c30c",
   18128 => x"30c30c",
   18129 => x"30c30c",
   18130 => x"30c30c",
   18131 => x"30c30c",
   18132 => x"30c30c",
   18133 => x"30c30c",
   18134 => x"30c30c",
   18135 => x"30c30c",
   18136 => x"30c30c",
   18137 => x"30c30c",
   18138 => x"30c30c",
   18139 => x"30c30c",
   18140 => x"30c30c",
   18141 => x"30c30c",
   18142 => x"30c30c",
   18143 => x"30c30c",
   18144 => x"30c30c",
   18145 => x"30c30c",
   18146 => x"30c30c",
   18147 => x"30c30c",
   18148 => x"77ffff",
   18149 => x"ffffff",
   18150 => x"ffffff",
   18151 => x"ffffff",
   18152 => x"ffffff",
   18153 => x"ffffff",
   18154 => x"ffffff",
   18155 => x"ffffff",
   18156 => x"ffffff",
   18157 => x"ffffff",
   18158 => x"ffffff",
   18159 => x"ffffff",
   18160 => x"ffffff",
   18161 => x"ffffff",
   18162 => x"ffffff",
   18163 => x"fea56a",
   18164 => x"ffffff",
   18165 => x"ffffff",
   18166 => x"ffffff",
   18167 => x"ffffff",
   18168 => x"ffffff",
   18169 => x"ffffff",
   18170 => x"ffffff",
   18171 => x"ffffff",
   18172 => x"ffffff",
   18173 => x"ffffff",
   18174 => x"ffffff",
   18175 => x"ffffff",
   18176 => x"ffffff",
   18177 => x"ffffff",
   18178 => x"ffffff",
   18179 => x"ffffff",
   18180 => x"ffffff",
   18181 => x"ffffff",
   18182 => x"ffffff",
   18183 => x"ffffff",
   18184 => x"ffffff",
   18185 => x"ffffff",
   18186 => x"ffffff",
   18187 => x"ffffff",
   18188 => x"ffffff",
   18189 => x"ffffff",
   18190 => x"ffffff",
   18191 => x"ffffff",
   18192 => x"ffffff",
   18193 => x"ffffff",
   18194 => x"ffffff",
   18195 => x"ffffff",
   18196 => x"ffffff",
   18197 => x"ffffff",
   18198 => x"ffffff",
   18199 => x"ffffff",
   18200 => x"ffffff",
   18201 => x"ffffff",
   18202 => x"ffffff",
   18203 => x"ffffff",
   18204 => x"ffffff",
   18205 => x"ffffff",
   18206 => x"ffffff",
   18207 => x"ffffff",
   18208 => x"ffffff",
   18209 => x"ffffff",
   18210 => x"ffffff",
   18211 => x"ffffff",
   18212 => x"ffffff",
   18213 => x"ffffff",
   18214 => x"ffffff",
   18215 => x"ffffff",
   18216 => x"ffffff",
   18217 => x"ffffff",
   18218 => x"ffffff",
   18219 => x"ffffff",
   18220 => x"ffffff",
   18221 => x"ffffff",
   18222 => x"ffffff",
   18223 => x"ffffff",
   18224 => x"ffffff",
   18225 => x"ffffff",
   18226 => x"ffffff",
   18227 => x"ffffff",
   18228 => x"ffffff",
   18229 => x"ffffff",
   18230 => x"ffffff",
   18231 => x"ffffff",
   18232 => x"ffffff",
   18233 => x"ffffff",
   18234 => x"ffffff",
   18235 => x"ffffff",
   18236 => x"ffffff",
   18237 => x"ffffff",
   18238 => x"ffffff",
   18239 => x"ffffff",
   18240 => x"ffac30",
   18241 => x"c30c30",
   18242 => x"c30c30",
   18243 => x"c30c30",
   18244 => x"c30c30",
   18245 => x"c30c30",
   18246 => x"c30c30",
   18247 => x"c30c30",
   18248 => x"c30c30",
   18249 => x"c30c30",
   18250 => x"c30c30",
   18251 => x"c30c30",
   18252 => x"c30c30",
   18253 => x"c30c30",
   18254 => x"c30c30",
   18255 => x"c30c30",
   18256 => x"c30c30",
   18257 => x"c30c30",
   18258 => x"c30c30",
   18259 => x"c30c30",
   18260 => x"c30c30",
   18261 => x"c30866",
   18262 => x"1abfff",
   18263 => x"ffffff",
   18264 => x"ffffff",
   18265 => x"ffffff",
   18266 => x"ffffff",
   18267 => x"ffffff",
   18268 => x"ffffff",
   18269 => x"ffffff",
   18270 => x"ffffff",
   18271 => x"ffffff",
   18272 => x"ffffff",
   18273 => x"ffffff",
   18274 => x"ffffff",
   18275 => x"ffffff",
   18276 => x"ffffff",
   18277 => x"ffffff",
   18278 => x"ffffff",
   18279 => x"ffffff",
   18280 => x"ffffff",
   18281 => x"ffffff",
   18282 => x"ffffff",
   18283 => x"ffffff",
   18284 => x"ffffff",
   18285 => x"ffffff",
   18286 => x"b8c38d",
   18287 => x"30c30c",
   18288 => x"30c30c",
   18289 => x"30c30c",
   18290 => x"30c30c",
   18291 => x"30c30c",
   18292 => x"30c30c",
   18293 => x"30c30c",
   18294 => x"30c30c",
   18295 => x"30c30c",
   18296 => x"30c30c",
   18297 => x"30c30c",
   18298 => x"30c30c",
   18299 => x"30c30c",
   18300 => x"30c30c",
   18301 => x"30c30c",
   18302 => x"30c30c",
   18303 => x"30c30c",
   18304 => x"30c30c",
   18305 => x"30c30c",
   18306 => x"30c30c",
   18307 => x"30c30c",
   18308 => x"77ffff",
   18309 => x"ffffff",
   18310 => x"ffffff",
   18311 => x"ffffff",
   18312 => x"ffffff",
   18313 => x"ffffff",
   18314 => x"ffffff",
   18315 => x"ffffff",
   18316 => x"ffffff",
   18317 => x"ffffff",
   18318 => x"ffffff",
   18319 => x"ffffff",
   18320 => x"ffffff",
   18321 => x"ffffff",
   18322 => x"ffffff",
   18323 => x"a95abf",
   18324 => x"ffffff",
   18325 => x"ffffff",
   18326 => x"ffffff",
   18327 => x"ffffff",
   18328 => x"ffffff",
   18329 => x"ffffff",
   18330 => x"ffffff",
   18331 => x"ffffff",
   18332 => x"ffffff",
   18333 => x"ffffff",
   18334 => x"ffffff",
   18335 => x"ffffff",
   18336 => x"ffffff",
   18337 => x"ffffff",
   18338 => x"ffffff",
   18339 => x"ffffff",
   18340 => x"ffffff",
   18341 => x"ffffff",
   18342 => x"ffffff",
   18343 => x"ffffff",
   18344 => x"ffffff",
   18345 => x"ffffff",
   18346 => x"ffffff",
   18347 => x"ffffff",
   18348 => x"ffffff",
   18349 => x"ffffff",
   18350 => x"ffffff",
   18351 => x"ffffff",
   18352 => x"ffffff",
   18353 => x"ffffff",
   18354 => x"ffffff",
   18355 => x"ffffff",
   18356 => x"ffffff",
   18357 => x"ffffff",
   18358 => x"ffffff",
   18359 => x"ffffff",
   18360 => x"ffffff",
   18361 => x"ffffff",
   18362 => x"ffffff",
   18363 => x"ffffff",
   18364 => x"ffffff",
   18365 => x"ffffff",
   18366 => x"ffffff",
   18367 => x"ffffff",
   18368 => x"ffffff",
   18369 => x"ffffff",
   18370 => x"ffffff",
   18371 => x"ffffff",
   18372 => x"ffffff",
   18373 => x"ffffff",
   18374 => x"ffffff",
   18375 => x"ffffff",
   18376 => x"ffffff",
   18377 => x"ffffff",
   18378 => x"ffffff",
   18379 => x"ffffff",
   18380 => x"ffffff",
   18381 => x"ffffff",
   18382 => x"ffffff",
   18383 => x"ffffff",
   18384 => x"ffffff",
   18385 => x"ffffff",
   18386 => x"ffffff",
   18387 => x"ffffff",
   18388 => x"ffffff",
   18389 => x"ffffff",
   18390 => x"ffffff",
   18391 => x"ffffff",
   18392 => x"ffffff",
   18393 => x"ffffff",
   18394 => x"ffffff",
   18395 => x"ffffff",
   18396 => x"ffffff",
   18397 => x"ffffff",
   18398 => x"ffffff",
   18399 => x"ffffff",
   18400 => x"fffc30",
   18401 => x"c30c30",
   18402 => x"c30c30",
   18403 => x"c30c30",
   18404 => x"c30c30",
   18405 => x"c30c30",
   18406 => x"c30c30",
   18407 => x"c30c30",
   18408 => x"c30c30",
   18409 => x"c30c30",
   18410 => x"c30c30",
   18411 => x"c30c30",
   18412 => x"c30c30",
   18413 => x"c30c30",
   18414 => x"c30c30",
   18415 => x"c30c30",
   18416 => x"c30c30",
   18417 => x"c30c30",
   18418 => x"c30c30",
   18419 => x"c30c30",
   18420 => x"c30c30",
   18421 => x"866aeb",
   18422 => x"5ebfff",
   18423 => x"ffffff",
   18424 => x"ffffff",
   18425 => x"ffffff",
   18426 => x"ffffff",
   18427 => x"ffffff",
   18428 => x"ffffff",
   18429 => x"ffffff",
   18430 => x"ffffff",
   18431 => x"ffffff",
   18432 => x"ffffff",
   18433 => x"ffffff",
   18434 => x"ffffff",
   18435 => x"ffffff",
   18436 => x"ffffff",
   18437 => x"ffffff",
   18438 => x"ffffff",
   18439 => x"ffffff",
   18440 => x"ffffff",
   18441 => x"ffffff",
   18442 => x"ffffff",
   18443 => x"ffffff",
   18444 => x"ffffff",
   18445 => x"ffffff",
   18446 => x"bcd3cf",
   18447 => x"38c30c",
   18448 => x"30c30c",
   18449 => x"30c30c",
   18450 => x"30c30c",
   18451 => x"30c30c",
   18452 => x"30c30c",
   18453 => x"30c30c",
   18454 => x"30c30c",
   18455 => x"30c30c",
   18456 => x"30c30c",
   18457 => x"30c30c",
   18458 => x"30c30c",
   18459 => x"30c30c",
   18460 => x"30c30c",
   18461 => x"30c30c",
   18462 => x"30c30c",
   18463 => x"30c30c",
   18464 => x"30c30c",
   18465 => x"30c30c",
   18466 => x"30c30c",
   18467 => x"30c30c",
   18468 => x"77ffff",
   18469 => x"ffffff",
   18470 => x"ffffff",
   18471 => x"ffffff",
   18472 => x"ffffff",
   18473 => x"ffffff",
   18474 => x"ffffff",
   18475 => x"ffffff",
   18476 => x"ffffff",
   18477 => x"ffffff",
   18478 => x"ffffff",
   18479 => x"ffffff",
   18480 => x"ffffff",
   18481 => x"ffffff",
   18482 => x"ffffea",
   18483 => x"56afff",
   18484 => x"ffffff",
   18485 => x"ffffff",
   18486 => x"ffffff",
   18487 => x"ffffff",
   18488 => x"ffffff",
   18489 => x"ffffff",
   18490 => x"ffffff",
   18491 => x"ffffff",
   18492 => x"ffffff",
   18493 => x"ffffff",
   18494 => x"ffffff",
   18495 => x"ffffff",
   18496 => x"ffffff",
   18497 => x"ffffff",
   18498 => x"ffffff",
   18499 => x"ffffff",
   18500 => x"ffffff",
   18501 => x"ffffff",
   18502 => x"ffffff",
   18503 => x"ffffff",
   18504 => x"ffffff",
   18505 => x"ffffff",
   18506 => x"ffffff",
   18507 => x"ffffff",
   18508 => x"ffffff",
   18509 => x"ffffff",
   18510 => x"ffffff",
   18511 => x"ffffff",
   18512 => x"ffffff",
   18513 => x"ffffff",
   18514 => x"ffffff",
   18515 => x"ffffff",
   18516 => x"ffffff",
   18517 => x"ffffff",
   18518 => x"ffffff",
   18519 => x"ffffff",
   18520 => x"ffffff",
   18521 => x"ffffff",
   18522 => x"ffffff",
   18523 => x"ffffff",
   18524 => x"ffffff",
   18525 => x"ffffff",
   18526 => x"ffffff",
   18527 => x"ffffff",
   18528 => x"ffffff",
   18529 => x"ffffff",
   18530 => x"ffffff",
   18531 => x"ffffff",
   18532 => x"ffffff",
   18533 => x"ffffff",
   18534 => x"ffffff",
   18535 => x"ffffff",
   18536 => x"ffffff",
   18537 => x"ffffff",
   18538 => x"ffffff",
   18539 => x"ffffff",
   18540 => x"ffffff",
   18541 => x"ffffff",
   18542 => x"ffffff",
   18543 => x"ffffff",
   18544 => x"ffffff",
   18545 => x"ffffff",
   18546 => x"ffffff",
   18547 => x"ffffff",
   18548 => x"ffffff",
   18549 => x"ffffff",
   18550 => x"ffffff",
   18551 => x"ffffff",
   18552 => x"ffffff",
   18553 => x"ffffff",
   18554 => x"ffffff",
   18555 => x"ffffff",
   18556 => x"ffffff",
   18557 => x"ffffff",
   18558 => x"ffffff",
   18559 => x"ffffff",
   18560 => x"fffc30",
   18561 => x"c30c30",
   18562 => x"c30c30",
   18563 => x"c30c30",
   18564 => x"c30c30",
   18565 => x"c30c30",
   18566 => x"c30c30",
   18567 => x"c30c30",
   18568 => x"c30c30",
   18569 => x"c30c30",
   18570 => x"c30c30",
   18571 => x"c30c30",
   18572 => x"c30c30",
   18573 => x"c30c30",
   18574 => x"c30c30",
   18575 => x"c30c30",
   18576 => x"c30c30",
   18577 => x"c30c30",
   18578 => x"c30c30",
   18579 => x"c30c30",
   18580 => x"c30c21",
   18581 => x"9a7df7",
   18582 => x"9eafff",
   18583 => x"ffffff",
   18584 => x"ffffff",
   18585 => x"ffffff",
   18586 => x"ffffff",
   18587 => x"ffffff",
   18588 => x"ffffff",
   18589 => x"ffffff",
   18590 => x"ffffff",
   18591 => x"ffffff",
   18592 => x"ffffff",
   18593 => x"ffffff",
   18594 => x"ffffff",
   18595 => x"ffffff",
   18596 => x"ffffff",
   18597 => x"ffffff",
   18598 => x"ffffff",
   18599 => x"ffffff",
   18600 => x"ffffff",
   18601 => x"ffffff",
   18602 => x"ffffff",
   18603 => x"ffffff",
   18604 => x"ffffff",
   18605 => x"ffffff",
   18606 => x"bcd3cf",
   18607 => x"3ce34c",
   18608 => x"30c30c",
   18609 => x"30c30c",
   18610 => x"30c30c",
   18611 => x"30c30c",
   18612 => x"30c30c",
   18613 => x"30c30c",
   18614 => x"30c30c",
   18615 => x"30c30c",
   18616 => x"30c30c",
   18617 => x"30c30c",
   18618 => x"30c30c",
   18619 => x"30c30c",
   18620 => x"30c30c",
   18621 => x"30c30c",
   18622 => x"30c30c",
   18623 => x"30c30c",
   18624 => x"30c30c",
   18625 => x"30c30c",
   18626 => x"30c30c",
   18627 => x"30c30c",
   18628 => x"bbffff",
   18629 => x"ffffff",
   18630 => x"ffffff",
   18631 => x"ffffff",
   18632 => x"ffffff",
   18633 => x"ffffff",
   18634 => x"ffffff",
   18635 => x"ffffff",
   18636 => x"ffffff",
   18637 => x"ffffff",
   18638 => x"ffffff",
   18639 => x"ffffff",
   18640 => x"ffffff",
   18641 => x"ffffff",
   18642 => x"fffa95",
   18643 => x"abffff",
   18644 => x"ffffff",
   18645 => x"ffffff",
   18646 => x"ffffff",
   18647 => x"ffffff",
   18648 => x"ffffff",
   18649 => x"ffffff",
   18650 => x"ffffff",
   18651 => x"ffffff",
   18652 => x"ffffff",
   18653 => x"ffffff",
   18654 => x"ffffff",
   18655 => x"ffffff",
   18656 => x"ffffff",
   18657 => x"ffffff",
   18658 => x"ffffff",
   18659 => x"ffffff",
   18660 => x"ffffff",
   18661 => x"ffffff",
   18662 => x"ffffff",
   18663 => x"ffffff",
   18664 => x"ffffff",
   18665 => x"ffffff",
   18666 => x"ffffff",
   18667 => x"ffffff",
   18668 => x"ffffff",
   18669 => x"ffffff",
   18670 => x"ffffff",
   18671 => x"ffffff",
   18672 => x"ffffff",
   18673 => x"ffffff",
   18674 => x"ffffff",
   18675 => x"ffffff",
   18676 => x"ffffff",
   18677 => x"ffffff",
   18678 => x"ffffff",
   18679 => x"ffffff",
   18680 => x"ffffff",
   18681 => x"ffffff",
   18682 => x"ffffff",
   18683 => x"ffffff",
   18684 => x"ffffff",
   18685 => x"ffffff",
   18686 => x"ffffff",
   18687 => x"ffffff",
   18688 => x"ffffff",
   18689 => x"ffffff",
   18690 => x"ffffff",
   18691 => x"ffffff",
   18692 => x"ffffff",
   18693 => x"ffffff",
   18694 => x"ffffff",
   18695 => x"ffffff",
   18696 => x"ffffff",
   18697 => x"ffffff",
   18698 => x"ffffff",
   18699 => x"ffffff",
   18700 => x"ffffff",
   18701 => x"ffffff",
   18702 => x"ffffff",
   18703 => x"ffffff",
   18704 => x"ffffff",
   18705 => x"ffffff",
   18706 => x"ffffff",
   18707 => x"ffffff",
   18708 => x"ffffff",
   18709 => x"ffffff",
   18710 => x"ffffff",
   18711 => x"ffffff",
   18712 => x"ffffff",
   18713 => x"ffffff",
   18714 => x"ffffff",
   18715 => x"ffffff",
   18716 => x"ffffff",
   18717 => x"ffffff",
   18718 => x"ffffff",
   18719 => x"ffffff",
   18720 => x"fffd70",
   18721 => x"c30c30",
   18722 => x"c30c30",
   18723 => x"c30c30",
   18724 => x"c30c30",
   18725 => x"c30c30",
   18726 => x"c30c30",
   18727 => x"c30c30",
   18728 => x"c30c30",
   18729 => x"c30c30",
   18730 => x"c30c30",
   18731 => x"c30c30",
   18732 => x"c30c30",
   18733 => x"c30c30",
   18734 => x"c30c30",
   18735 => x"c30c30",
   18736 => x"c30c30",
   18737 => x"c30c30",
   18738 => x"c30c30",
   18739 => x"c30c30",
   18740 => x"c309a7",
   18741 => x"df3cf3",
   18742 => x"9dabbf",
   18743 => x"ffffff",
   18744 => x"ffffff",
   18745 => x"ffffff",
   18746 => x"ffffff",
   18747 => x"ffffff",
   18748 => x"ffffff",
   18749 => x"ffffff",
   18750 => x"ffffff",
   18751 => x"ffffff",
   18752 => x"ffffff",
   18753 => x"ffffff",
   18754 => x"ffffff",
   18755 => x"ffffff",
   18756 => x"ffffff",
   18757 => x"ffffff",
   18758 => x"ffffff",
   18759 => x"ffffff",
   18760 => x"ffffff",
   18761 => x"ffffff",
   18762 => x"ffffff",
   18763 => x"ffffff",
   18764 => x"ffffff",
   18765 => x"ffffff",
   18766 => x"b8e3cf",
   18767 => x"3cf38d",
   18768 => x"30c30c",
   18769 => x"30c30c",
   18770 => x"30c30c",
   18771 => x"30c30c",
   18772 => x"30c30c",
   18773 => x"30c30c",
   18774 => x"30c30c",
   18775 => x"30c30c",
   18776 => x"30c30c",
   18777 => x"30c30c",
   18778 => x"30c30c",
   18779 => x"30c30c",
   18780 => x"30c30c",
   18781 => x"30c30c",
   18782 => x"30c30c",
   18783 => x"30c30c",
   18784 => x"30c30c",
   18785 => x"30c30c",
   18786 => x"30c30c",
   18787 => x"30c30c",
   18788 => x"bbffff",
   18789 => x"ffffff",
   18790 => x"ffffff",
   18791 => x"ffffff",
   18792 => x"ffffff",
   18793 => x"ffffff",
   18794 => x"ffffff",
   18795 => x"ffffff",
   18796 => x"ffffff",
   18797 => x"ffffff",
   18798 => x"ffffff",
   18799 => x"ffffff",
   18800 => x"ffffff",
   18801 => x"ffffff",
   18802 => x"fea56a",
   18803 => x"ffffff",
   18804 => x"ffffff",
   18805 => x"ffffff",
   18806 => x"ffffff",
   18807 => x"ffffff",
   18808 => x"ffffff",
   18809 => x"ffffff",
   18810 => x"ffffff",
   18811 => x"ffffff",
   18812 => x"ffffff",
   18813 => x"ffffff",
   18814 => x"ffffff",
   18815 => x"ffffff",
   18816 => x"ffffff",
   18817 => x"ffffff",
   18818 => x"ffffff",
   18819 => x"ffffff",
   18820 => x"ffffff",
   18821 => x"ffffff",
   18822 => x"ffffff",
   18823 => x"ffffff",
   18824 => x"ffffff",
   18825 => x"ffffff",
   18826 => x"ffffff",
   18827 => x"ffffff",
   18828 => x"ffffff",
   18829 => x"ffffff",
   18830 => x"ffffff",
   18831 => x"ffffff",
   18832 => x"ffffff",
   18833 => x"ffffff",
   18834 => x"ffffff",
   18835 => x"ffffff",
   18836 => x"ffffff",
   18837 => x"ffffff",
   18838 => x"ffffff",
   18839 => x"ffffff",
   18840 => x"ffffff",
   18841 => x"ffffff",
   18842 => x"ffffff",
   18843 => x"ffffff",
   18844 => x"ffffff",
   18845 => x"ffffff",
   18846 => x"ffffff",
   18847 => x"ffffff",
   18848 => x"ffffff",
   18849 => x"ffffff",
   18850 => x"ffffff",
   18851 => x"ffffff",
   18852 => x"ffffff",
   18853 => x"ffffff",
   18854 => x"ffffff",
   18855 => x"ffffff",
   18856 => x"ffffff",
   18857 => x"ffffff",
   18858 => x"ffffff",
   18859 => x"ffffff",
   18860 => x"ffffff",
   18861 => x"ffffff",
   18862 => x"ffffff",
   18863 => x"ffffff",
   18864 => x"ffffff",
   18865 => x"ffffff",
   18866 => x"ffffff",
   18867 => x"ffffff",
   18868 => x"ffffff",
   18869 => x"ffffff",
   18870 => x"ffffff",
   18871 => x"ffffff",
   18872 => x"ffffff",
   18873 => x"ffffff",
   18874 => x"ffffff",
   18875 => x"ffffff",
   18876 => x"ffffff",
   18877 => x"ffffff",
   18878 => x"ffffff",
   18879 => x"ffffff",
   18880 => x"fffd70",
   18881 => x"c30c30",
   18882 => x"c30c30",
   18883 => x"c30c30",
   18884 => x"c30c30",
   18885 => x"c30c30",
   18886 => x"c30c30",
   18887 => x"c30c30",
   18888 => x"c30c30",
   18889 => x"c30c30",
   18890 => x"c30c30",
   18891 => x"c30c30",
   18892 => x"c30c30",
   18893 => x"c30c30",
   18894 => x"c30c30",
   18895 => x"c30c30",
   18896 => x"c30c30",
   18897 => x"c30c30",
   18898 => x"c30c30",
   18899 => x"c30c30",
   18900 => x"8669f7",
   18901 => x"cf3cf3",
   18902 => x"ddabbf",
   18903 => x"ffffff",
   18904 => x"ffffff",
   18905 => x"ffffff",
   18906 => x"ffffff",
   18907 => x"ffffff",
   18908 => x"ffffff",
   18909 => x"ffffff",
   18910 => x"ffffff",
   18911 => x"ffffff",
   18912 => x"ffffff",
   18913 => x"ffffff",
   18914 => x"ffffff",
   18915 => x"ffffff",
   18916 => x"ffffff",
   18917 => x"ffffff",
   18918 => x"ffffff",
   18919 => x"ffffff",
   18920 => x"ffffff",
   18921 => x"ffffff",
   18922 => x"ffffff",
   18923 => x"ffffff",
   18924 => x"ffffff",
   18925 => x"ffffff",
   18926 => x"b8e3cf",
   18927 => x"3cf3cf",
   18928 => x"38c30c",
   18929 => x"30c30c",
   18930 => x"30c30c",
   18931 => x"30c30c",
   18932 => x"30c30c",
   18933 => x"30c30c",
   18934 => x"30c30c",
   18935 => x"30c30c",
   18936 => x"30c30c",
   18937 => x"30c30c",
   18938 => x"30c30c",
   18939 => x"30c30c",
   18940 => x"30c30c",
   18941 => x"30c30c",
   18942 => x"30c30c",
   18943 => x"30c30c",
   18944 => x"30c30c",
   18945 => x"30c30c",
   18946 => x"30c30c",
   18947 => x"30c30c",
   18948 => x"bbffff",
   18949 => x"ffffff",
   18950 => x"ffffff",
   18951 => x"ffffff",
   18952 => x"ffffff",
   18953 => x"ffffff",
   18954 => x"ffffff",
   18955 => x"ffffff",
   18956 => x"ffffff",
   18957 => x"ffffff",
   18958 => x"ffffff",
   18959 => x"ffffff",
   18960 => x"ffffff",
   18961 => x"ffffff",
   18962 => x"a95abf",
   18963 => x"ffffff",
   18964 => x"ffffff",
   18965 => x"ffffff",
   18966 => x"ffffff",
   18967 => x"ffffff",
   18968 => x"ffffff",
   18969 => x"ffffff",
   18970 => x"ffffff",
   18971 => x"ffffff",
   18972 => x"ffffff",
   18973 => x"ffffff",
   18974 => x"ffffff",
   18975 => x"ffffff",
   18976 => x"ffffff",
   18977 => x"ffffff",
   18978 => x"ffffff",
   18979 => x"ffffff",
   18980 => x"ffffff",
   18981 => x"ffffff",
   18982 => x"ffffff",
   18983 => x"ffffff",
   18984 => x"ffffff",
   18985 => x"ffffff",
   18986 => x"ffffff",
   18987 => x"ffffff",
   18988 => x"ffffff",
   18989 => x"ffffff",
   18990 => x"ffffff",
   18991 => x"ffffff",
   18992 => x"ffffff",
   18993 => x"ffffff",
   18994 => x"ffffff",
   18995 => x"ffffff",
   18996 => x"ffffff",
   18997 => x"ffffff",
   18998 => x"ffffff",
   18999 => x"ffffff",
   19000 => x"ffffff",
   19001 => x"ffffff",
   19002 => x"ffffff",
   19003 => x"ffffff",
   19004 => x"ffffff",
   19005 => x"ffffff",
   19006 => x"ffffff",
   19007 => x"ffffff",
   19008 => x"ffffff",
   19009 => x"ffffff",
   19010 => x"ffffff",
   19011 => x"ffffff",
   19012 => x"ffffff",
   19013 => x"ffffff",
   19014 => x"ffffff",
   19015 => x"ffffff",
   19016 => x"ffffff",
   19017 => x"ffffff",
   19018 => x"ffffff",
   19019 => x"ffffff",
   19020 => x"ffffff",
   19021 => x"ffffff",
   19022 => x"ffffff",
   19023 => x"ffffff",
   19024 => x"ffffff",
   19025 => x"ffffff",
   19026 => x"ffffff",
   19027 => x"ffffff",
   19028 => x"ffffff",
   19029 => x"ffffff",
   19030 => x"ffffff",
   19031 => x"ffffff",
   19032 => x"ffffff",
   19033 => x"ffffff",
   19034 => x"ffffff",
   19035 => x"ffffff",
   19036 => x"ffffff",
   19037 => x"ffffff",
   19038 => x"ffffff",
   19039 => x"ffffff",
   19040 => x"fffeb0",
   19041 => x"c30c30",
   19042 => x"c30c30",
   19043 => x"c30c30",
   19044 => x"c30c30",
   19045 => x"c30c30",
   19046 => x"c30c30",
   19047 => x"c30c30",
   19048 => x"c30c30",
   19049 => x"c30c30",
   19050 => x"c30c30",
   19051 => x"c30c30",
   19052 => x"c30c30",
   19053 => x"c30c30",
   19054 => x"c30c30",
   19055 => x"c30c30",
   19056 => x"c30c30",
   19057 => x"c30c30",
   19058 => x"c30c30",
   19059 => x"c30c21",
   19060 => x"9a7cf3",
   19061 => x"cf3cf3",
   19062 => x"ddabbf",
   19063 => x"ffffff",
   19064 => x"ffffff",
   19065 => x"ffffff",
   19066 => x"ffffff",
   19067 => x"ffffff",
   19068 => x"ffffff",
   19069 => x"ffffff",
   19070 => x"ffffff",
   19071 => x"ffffff",
   19072 => x"ffffff",
   19073 => x"ffffff",
   19074 => x"ffffff",
   19075 => x"ffffff",
   19076 => x"ffffff",
   19077 => x"ffffff",
   19078 => x"ffffff",
   19079 => x"ffffff",
   19080 => x"ffffff",
   19081 => x"ffffff",
   19082 => x"ffffff",
   19083 => x"ffffff",
   19084 => x"ffffff",
   19085 => x"ffffff",
   19086 => x"78f3cf",
   19087 => x"3cf3cf",
   19088 => x"3ce34c",
   19089 => x"30c30c",
   19090 => x"30c30c",
   19091 => x"30c30c",
   19092 => x"30c30c",
   19093 => x"30c30c",
   19094 => x"30c30c",
   19095 => x"30c30c",
   19096 => x"30c30c",
   19097 => x"30c30c",
   19098 => x"30c30c",
   19099 => x"30c30c",
   19100 => x"30c30c",
   19101 => x"30c30c",
   19102 => x"30c30c",
   19103 => x"30c30c",
   19104 => x"30c30c",
   19105 => x"30c30c",
   19106 => x"30c30c",
   19107 => x"30c30c",
   19108 => x"bbffff",
   19109 => x"ffffff",
   19110 => x"ffffff",
   19111 => x"ffffff",
   19112 => x"ffffff",
   19113 => x"ffffff",
   19114 => x"ffffff",
   19115 => x"ffffff",
   19116 => x"ffffff",
   19117 => x"ffffff",
   19118 => x"ffffff",
   19119 => x"ffffff",
   19120 => x"ffffff",
   19121 => x"ffffea",
   19122 => x"56afff",
   19123 => x"ffffff",
   19124 => x"ffffff",
   19125 => x"ffffff",
   19126 => x"ffffff",
   19127 => x"ffffff",
   19128 => x"ffffff",
   19129 => x"ffffff",
   19130 => x"ffffff",
   19131 => x"ffffff",
   19132 => x"ffffff",
   19133 => x"ffffff",
   19134 => x"ffffff",
   19135 => x"ffffff",
   19136 => x"ffffff",
   19137 => x"ffffff",
   19138 => x"ffffff",
   19139 => x"ffffff",
   19140 => x"ffffff",
   19141 => x"ffffff",
   19142 => x"ffffff",
   19143 => x"ffffff",
   19144 => x"ffffff",
   19145 => x"ffffff",
   19146 => x"ffffff",
   19147 => x"ffffff",
   19148 => x"ffffff",
   19149 => x"ffffff",
   19150 => x"ffffff",
   19151 => x"ffffff",
   19152 => x"ffffff",
   19153 => x"ffffff",
   19154 => x"ffffff",
   19155 => x"ffffff",
   19156 => x"ffffff",
   19157 => x"ffffff",
   19158 => x"ffffff",
   19159 => x"ffffff",
   19160 => x"ffffff",
   19161 => x"ffffff",
   19162 => x"ffffff",
   19163 => x"ffffff",
   19164 => x"ffffff",
   19165 => x"ffffff",
   19166 => x"ffffff",
   19167 => x"ffffff",
   19168 => x"ffffff",
   19169 => x"ffffff",
   19170 => x"ffffff",
   19171 => x"ffffff",
   19172 => x"ffffff",
   19173 => x"ffffff",
   19174 => x"ffffff",
   19175 => x"ffffff",
   19176 => x"ffffff",
   19177 => x"ffffff",
   19178 => x"ffffff",
   19179 => x"ffffff",
   19180 => x"ffffff",
   19181 => x"ffffff",
   19182 => x"ffffff",
   19183 => x"ffffff",
   19184 => x"ffffff",
   19185 => x"ffffff",
   19186 => x"ffffff",
   19187 => x"ffffff",
   19188 => x"ffffff",
   19189 => x"ffffff",
   19190 => x"ffffff",
   19191 => x"ffffff",
   19192 => x"ffffff",
   19193 => x"ffffff",
   19194 => x"ffffff",
   19195 => x"ffffff",
   19196 => x"ffffff",
   19197 => x"ffffff",
   19198 => x"ffffff",
   19199 => x"ffffff",
   19200 => x"fffeb0",
   19201 => x"c30c30",
   19202 => x"c30c30",
   19203 => x"c30c30",
   19204 => x"c30c30",
   19205 => x"c30c30",
   19206 => x"c30c30",
   19207 => x"c30c30",
   19208 => x"c30c30",
   19209 => x"c30c30",
   19210 => x"c30c30",
   19211 => x"c30c30",
   19212 => x"c30c30",
   19213 => x"c30c30",
   19214 => x"c30c30",
   19215 => x"c30c30",
   19216 => x"c30c30",
   19217 => x"c30c30",
   19218 => x"c30c30",
   19219 => x"c30867",
   19220 => x"df3cf3",
   19221 => x"cf3cf3",
   19222 => x"cd6bbf",
   19223 => x"ffffff",
   19224 => x"ffffff",
   19225 => x"ffffff",
   19226 => x"ffffff",
   19227 => x"ffffff",
   19228 => x"ffffff",
   19229 => x"ffffff",
   19230 => x"ffffff",
   19231 => x"ffffff",
   19232 => x"ffffff",
   19233 => x"ffffff",
   19234 => x"ffffff",
   19235 => x"ffffff",
   19236 => x"ffffff",
   19237 => x"ffffff",
   19238 => x"ffffff",
   19239 => x"ffffff",
   19240 => x"ffffff",
   19241 => x"ffffff",
   19242 => x"ffffff",
   19243 => x"ffffff",
   19244 => x"ffffff",
   19245 => x"ffffff",
   19246 => x"78f3cf",
   19247 => x"3cf3cf",
   19248 => x"3cf38d",
   19249 => x"30c30c",
   19250 => x"30c30c",
   19251 => x"30c30c",
   19252 => x"30c30c",
   19253 => x"30c30c",
   19254 => x"30c30c",
   19255 => x"30c30c",
   19256 => x"30c30c",
   19257 => x"30c30c",
   19258 => x"30c30c",
   19259 => x"30c30c",
   19260 => x"30c30c",
   19261 => x"30c30c",
   19262 => x"30c30c",
   19263 => x"30c30c",
   19264 => x"30c30c",
   19265 => x"30c30c",
   19266 => x"30c30c",
   19267 => x"30c31d",
   19268 => x"ffffff",
   19269 => x"ffffff",
   19270 => x"ffffff",
   19271 => x"ffffff",
   19272 => x"ffffff",
   19273 => x"ffffff",
   19274 => x"ffffff",
   19275 => x"ffffff",
   19276 => x"ffffff",
   19277 => x"ffffff",
   19278 => x"ffffff",
   19279 => x"ffffff",
   19280 => x"ffffff",
   19281 => x"fffa95",
   19282 => x"abffff",
   19283 => x"ffffff",
   19284 => x"ffffff",
   19285 => x"ffffff",
   19286 => x"ffffff",
   19287 => x"ffffff",
   19288 => x"ffffff",
   19289 => x"ffffff",
   19290 => x"ffffff",
   19291 => x"ffffff",
   19292 => x"ffffff",
   19293 => x"ffffff",
   19294 => x"ffffff",
   19295 => x"ffffff",
   19296 => x"ffffff",
   19297 => x"ffffff",
   19298 => x"ffffff",
   19299 => x"ffffff",
   19300 => x"ffffff",
   19301 => x"ffffff",
   19302 => x"ffffff",
   19303 => x"ffffff",
   19304 => x"ffffff",
   19305 => x"ffffff",
   19306 => x"ffffff",
   19307 => x"ffffff",
   19308 => x"ffffff",
   19309 => x"ffffff",
   19310 => x"ffffff",
   19311 => x"ffffff",
   19312 => x"ffffff",
   19313 => x"ffffff",
   19314 => x"ffffff",
   19315 => x"ffffff",
   19316 => x"ffffff",
   19317 => x"ffffff",
   19318 => x"ffffff",
   19319 => x"ffffff",
   19320 => x"ffffff",
   19321 => x"ffffff",
   19322 => x"ffffff",
   19323 => x"ffffff",
   19324 => x"ffffff",
   19325 => x"ffffff",
   19326 => x"ffffff",
   19327 => x"ffffff",
   19328 => x"ffffff",
   19329 => x"ffffff",
   19330 => x"ffffff",
   19331 => x"ffffff",
   19332 => x"ffffff",
   19333 => x"ffffff",
   19334 => x"ffffff",
   19335 => x"ffffff",
   19336 => x"ffffff",
   19337 => x"ffffff",
   19338 => x"ffffff",
   19339 => x"ffffff",
   19340 => x"ffffff",
   19341 => x"ffffff",
   19342 => x"ffffff",
   19343 => x"ffffff",
   19344 => x"ffffff",
   19345 => x"ffffff",
   19346 => x"ffffff",
   19347 => x"ffffff",
   19348 => x"ffffff",
   19349 => x"ffffff",
   19350 => x"ffffff",
   19351 => x"ffffff",
   19352 => x"ffffff",
   19353 => x"ffffff",
   19354 => x"ffffff",
   19355 => x"ffffff",
   19356 => x"ffffff",
   19357 => x"ffffff",
   19358 => x"ffffff",
   19359 => x"ffffff",
   19360 => x"fffeb0",
   19361 => x"c30c30",
   19362 => x"c30c30",
   19363 => x"c30c30",
   19364 => x"c30c30",
   19365 => x"c30c30",
   19366 => x"c30c30",
   19367 => x"c30c30",
   19368 => x"c30c30",
   19369 => x"c30c30",
   19370 => x"c30c30",
   19371 => x"c30c30",
   19372 => x"c30c30",
   19373 => x"c30c30",
   19374 => x"c30c30",
   19375 => x"c30c30",
   19376 => x"c30c30",
   19377 => x"c30c30",
   19378 => x"c30c30",
   19379 => x"c229f7",
   19380 => x"cf3cf3",
   19381 => x"cf3cf3",
   19382 => x"ce7bbf",
   19383 => x"ffffff",
   19384 => x"ffffff",
   19385 => x"ffffff",
   19386 => x"ffffff",
   19387 => x"ffffff",
   19388 => x"ffffff",
   19389 => x"ffffff",
   19390 => x"ffffff",
   19391 => x"ffffff",
   19392 => x"ffffff",
   19393 => x"ffffff",
   19394 => x"ffffff",
   19395 => x"ffffff",
   19396 => x"ffffff",
   19397 => x"ffffff",
   19398 => x"ffffff",
   19399 => x"ffffff",
   19400 => x"ffffff",
   19401 => x"ffffff",
   19402 => x"ffffff",
   19403 => x"ffffff",
   19404 => x"ffffff",
   19405 => x"ffffff",
   19406 => x"78f3cf",
   19407 => x"3cf3cf",
   19408 => x"3cf3ce",
   19409 => x"34c30c",
   19410 => x"30c30c",
   19411 => x"30c30c",
   19412 => x"30c30c",
   19413 => x"30c30c",
   19414 => x"30c30c",
   19415 => x"30c30c",
   19416 => x"30c30c",
   19417 => x"30c30c",
   19418 => x"30c30c",
   19419 => x"30c30c",
   19420 => x"30c30c",
   19421 => x"30c30c",
   19422 => x"30c30c",
   19423 => x"30c30c",
   19424 => x"30c30c",
   19425 => x"30c30c",
   19426 => x"30c30c",
   19427 => x"30c31d",
   19428 => x"ffffff",
   19429 => x"ffffff",
   19430 => x"ffffff",
   19431 => x"ffffff",
   19432 => x"ffffff",
   19433 => x"ffffff",
   19434 => x"ffffff",
   19435 => x"ffffff",
   19436 => x"ffffff",
   19437 => x"ffffff",
   19438 => x"ffffff",
   19439 => x"ffffff",
   19440 => x"ffffff",
   19441 => x"fea56a",
   19442 => x"ffffff",
   19443 => x"ffffff",
   19444 => x"ffffff",
   19445 => x"ffffff",
   19446 => x"ffffff",
   19447 => x"ffffff",
   19448 => x"ffffff",
   19449 => x"ffffff",
   19450 => x"ffffff",
   19451 => x"ffffff",
   19452 => x"ffffff",
   19453 => x"ffffff",
   19454 => x"ffffff",
   19455 => x"ffffff",
   19456 => x"ffffff",
   19457 => x"ffffff",
   19458 => x"ffffff",
   19459 => x"ffffff",
   19460 => x"ffffff",
   19461 => x"ffffff",
   19462 => x"ffffff",
   19463 => x"ffffff",
   19464 => x"ffffff",
   19465 => x"ffffff",
   19466 => x"ffffff",
   19467 => x"ffffff",
   19468 => x"ffffff",
   19469 => x"ffffff",
   19470 => x"ffffff",
   19471 => x"ffffff",
   19472 => x"ffffff",
   19473 => x"ffffff",
   19474 => x"ffffff",
   19475 => x"ffffff",
   19476 => x"ffffff",
   19477 => x"ffffff",
   19478 => x"ffffff",
   19479 => x"ffffff",
   19480 => x"ffffff",
   19481 => x"ffffff",
   19482 => x"ffffff",
   19483 => x"ffffff",
   19484 => x"ffffff",
   19485 => x"ffffff",
   19486 => x"ffffff",
   19487 => x"ffffff",
   19488 => x"ffffff",
   19489 => x"ffffff",
   19490 => x"ffffff",
   19491 => x"ffffff",
   19492 => x"ffffff",
   19493 => x"ffffff",
   19494 => x"ffffff",
   19495 => x"ffffff",
   19496 => x"ffffff",
   19497 => x"ffffff",
   19498 => x"ffffff",
   19499 => x"ffffff",
   19500 => x"ffffff",
   19501 => x"ffffff",
   19502 => x"ffffff",
   19503 => x"ffffff",
   19504 => x"ffffff",
   19505 => x"ffffff",
   19506 => x"ffffff",
   19507 => x"ffffff",
   19508 => x"ffffff",
   19509 => x"ffffff",
   19510 => x"ffffff",
   19511 => x"ffffff",
   19512 => x"ffffff",
   19513 => x"ffffff",
   19514 => x"ffffff",
   19515 => x"ffffff",
   19516 => x"ffffff",
   19517 => x"ffffff",
   19518 => x"ffffff",
   19519 => x"ffffff",
   19520 => x"fffff0",
   19521 => x"c30c30",
   19522 => x"c30c30",
   19523 => x"c30c30",
   19524 => x"c30c30",
   19525 => x"c30c30",
   19526 => x"c30c30",
   19527 => x"c30c30",
   19528 => x"c30c30",
   19529 => x"c30c30",
   19530 => x"c30c30",
   19531 => x"c30c30",
   19532 => x"c30c30",
   19533 => x"c30c30",
   19534 => x"c30c30",
   19535 => x"c30c30",
   19536 => x"c30c30",
   19537 => x"c30c30",
   19538 => x"c30c30",
   19539 => x"8a7df3",
   19540 => x"cf3cf3",
   19541 => x"cf3cf3",
   19542 => x"cf7aae",
   19543 => x"ffffff",
   19544 => x"ffffff",
   19545 => x"ffffff",
   19546 => x"ffffff",
   19547 => x"ffffff",
   19548 => x"ffffff",
   19549 => x"ffffff",
   19550 => x"ffffff",
   19551 => x"ffffff",
   19552 => x"ffffff",
   19553 => x"ffffff",
   19554 => x"ffffff",
   19555 => x"ffffff",
   19556 => x"ffffff",
   19557 => x"ffffff",
   19558 => x"ffffff",
   19559 => x"ffffff",
   19560 => x"ffffff",
   19561 => x"ffffff",
   19562 => x"ffffff",
   19563 => x"ffffff",
   19564 => x"ffffff",
   19565 => x"ffffef",
   19566 => x"38f3cf",
   19567 => x"3cf3cf",
   19568 => x"3cf3cf",
   19569 => x"3cd30c",
   19570 => x"30c30c",
   19571 => x"30c30c",
   19572 => x"30c30c",
   19573 => x"30c30c",
   19574 => x"30c30c",
   19575 => x"30c30c",
   19576 => x"30c30c",
   19577 => x"30c30c",
   19578 => x"30c30c",
   19579 => x"30c30c",
   19580 => x"30c30c",
   19581 => x"30c30c",
   19582 => x"30c30c",
   19583 => x"30c30c",
   19584 => x"30c30c",
   19585 => x"30c30c",
   19586 => x"30c30c",
   19587 => x"30c32e",
   19588 => x"ffffff",
   19589 => x"ffffff",
   19590 => x"ffffff",
   19591 => x"ffffff",
   19592 => x"ffffff",
   19593 => x"ffffff",
   19594 => x"ffffff",
   19595 => x"ffffff",
   19596 => x"ffffff",
   19597 => x"ffffff",
   19598 => x"ffffff",
   19599 => x"ffffff",
   19600 => x"ffffff",
   19601 => x"a95abf",
   19602 => x"ffffff",
   19603 => x"ffffff",
   19604 => x"ffffff",
   19605 => x"ffffff",
   19606 => x"ffffff",
   19607 => x"ffffff",
   19608 => x"ffffff",
   19609 => x"ffffff",
   19610 => x"ffffff",
   19611 => x"ffffff",
   19612 => x"ffffff",
   19613 => x"ffffff",
   19614 => x"ffffff",
   19615 => x"ffffff",
   19616 => x"ffffff",
   19617 => x"ffffff",
   19618 => x"ffffff",
   19619 => x"ffffff",
   19620 => x"ffffff",
   19621 => x"ffffff",
   19622 => x"ffffff",
   19623 => x"ffffff",
   19624 => x"ffffff",
   19625 => x"ffffff",
   19626 => x"ffffff",
   19627 => x"ffffff",
   19628 => x"ffffff",
   19629 => x"ffffff",
   19630 => x"ffffff",
   19631 => x"ffffff",
   19632 => x"ffffff",
   19633 => x"ffffff",
   19634 => x"ffffff",
   19635 => x"ffffff",
   19636 => x"ffffff",
   19637 => x"ffffff",
   19638 => x"ffffff",
   19639 => x"ffffff",
   19640 => x"ffffff",
   19641 => x"ffffff",
   19642 => x"ffffff",
   19643 => x"ffffff",
   19644 => x"ffffff",
   19645 => x"ffffff",
   19646 => x"ffffff",
   19647 => x"ffffff",
   19648 => x"ffffff",
   19649 => x"ffffff",
   19650 => x"ffffff",
   19651 => x"ffffff",
   19652 => x"ffffff",
   19653 => x"ffffff",
   19654 => x"ffffff",
   19655 => x"ffffff",
   19656 => x"ffffff",
   19657 => x"ffffff",
   19658 => x"ffffff",
   19659 => x"ffffff",
   19660 => x"ffffff",
   19661 => x"ffffff",
   19662 => x"ffffff",
   19663 => x"ffffff",
   19664 => x"ffffff",
   19665 => x"ffffff",
   19666 => x"ffffff",
   19667 => x"ffffff",
   19668 => x"ffffff",
   19669 => x"ffffff",
   19670 => x"ffffff",
   19671 => x"ffffff",
   19672 => x"ffffff",
   19673 => x"ffffff",
   19674 => x"ffffff",
   19675 => x"ffffff",
   19676 => x"ffffff",
   19677 => x"ffffff",
   19678 => x"ffffff",
   19679 => x"ffffff",
   19680 => x"fffff5",
   19681 => x"c30c30",
   19682 => x"c30c30",
   19683 => x"c30c30",
   19684 => x"c30c30",
   19685 => x"c30c30",
   19686 => x"c30c30",
   19687 => x"c30c30",
   19688 => x"c30c30",
   19689 => x"c30c30",
   19690 => x"c30c30",
   19691 => x"c30c30",
   19692 => x"c30c30",
   19693 => x"c30c30",
   19694 => x"c30c30",
   19695 => x"c30c30",
   19696 => x"c30c30",
   19697 => x"c30c30",
   19698 => x"c30866",
   19699 => x"9f7cf3",
   19700 => x"cf3cf3",
   19701 => x"cf3cf3",
   19702 => x"cf7aae",
   19703 => x"ffffff",
   19704 => x"ffffff",
   19705 => x"ffffff",
   19706 => x"ffffff",
   19707 => x"ffffff",
   19708 => x"ffffff",
   19709 => x"ffffff",
   19710 => x"ffffff",
   19711 => x"ffffff",
   19712 => x"ffffff",
   19713 => x"ffffff",
   19714 => x"ffffff",
   19715 => x"ffffff",
   19716 => x"ffffff",
   19717 => x"ffffff",
   19718 => x"ffffff",
   19719 => x"ffffff",
   19720 => x"ffffff",
   19721 => x"ffffff",
   19722 => x"ffffff",
   19723 => x"ffffff",
   19724 => x"ffffff",
   19725 => x"ffffee",
   19726 => x"38f3cf",
   19727 => x"3cf3cf",
   19728 => x"3cf3cf",
   19729 => x"3cf38c",
   19730 => x"30c30c",
   19731 => x"30c30c",
   19732 => x"30c30c",
   19733 => x"30c30c",
   19734 => x"30c30c",
   19735 => x"30c30c",
   19736 => x"30c30c",
   19737 => x"30c30c",
   19738 => x"30c30c",
   19739 => x"30c30c",
   19740 => x"30c30c",
   19741 => x"30c30c",
   19742 => x"30c30c",
   19743 => x"30c30c",
   19744 => x"30c30c",
   19745 => x"30c30c",
   19746 => x"30c30c",
   19747 => x"30c32e",
   19748 => x"ffffff",
   19749 => x"ffffff",
   19750 => x"ffffff",
   19751 => x"ffffff",
   19752 => x"ffffff",
   19753 => x"ffffff",
   19754 => x"ffffff",
   19755 => x"ffffff",
   19756 => x"ffffff",
   19757 => x"ffffff",
   19758 => x"ffffff",
   19759 => x"ffffff",
   19760 => x"ffffea",
   19761 => x"56afff",
   19762 => x"ffffff",
   19763 => x"ffffff",
   19764 => x"ffffff",
   19765 => x"ffffff",
   19766 => x"ffffff",
   19767 => x"ffffff",
   19768 => x"ffffff",
   19769 => x"ffffff",
   19770 => x"ffffff",
   19771 => x"ffffff",
   19772 => x"ffffff",
   19773 => x"ffffff",
   19774 => x"ffffff",
   19775 => x"ffffff",
   19776 => x"ffffff",
   19777 => x"ffffff",
   19778 => x"ffffff",
   19779 => x"ffffff",
   19780 => x"ffffff",
   19781 => x"ffffff",
   19782 => x"ffffff",
   19783 => x"ffffff",
   19784 => x"ffffff",
   19785 => x"ffffff",
   19786 => x"ffffff",
   19787 => x"ffffff",
   19788 => x"ffffff",
   19789 => x"ffffff",
   19790 => x"ffffff",
   19791 => x"ffffff",
   19792 => x"ffffff",
   19793 => x"ffffff",
   19794 => x"ffffff",
   19795 => x"ffffff",
   19796 => x"ffffff",
   19797 => x"ffffff",
   19798 => x"ffffff",
   19799 => x"ffffff",
   19800 => x"ffffff",
   19801 => x"ffffff",
   19802 => x"ffffff",
   19803 => x"ffffff",
   19804 => x"ffffff",
   19805 => x"ffffff",
   19806 => x"ffffff",
   19807 => x"ffffff",
   19808 => x"ffffff",
   19809 => x"ffffff",
   19810 => x"ffffff",
   19811 => x"ffffff",
   19812 => x"ffffff",
   19813 => x"ffffff",
   19814 => x"ffffff",
   19815 => x"ffffff",
   19816 => x"ffffff",
   19817 => x"ffffff",
   19818 => x"ffffff",
   19819 => x"ffffff",
   19820 => x"ffffff",
   19821 => x"ffffff",
   19822 => x"ffffff",
   19823 => x"ffffff",
   19824 => x"ffffff",
   19825 => x"ffffff",
   19826 => x"ffffff",
   19827 => x"ffffff",
   19828 => x"ffffff",
   19829 => x"ffffff",
   19830 => x"ffffff",
   19831 => x"ffffff",
   19832 => x"ffffff",
   19833 => x"ffffff",
   19834 => x"ffffff",
   19835 => x"ffffff",
   19836 => x"ffffff",
   19837 => x"ffffff",
   19838 => x"ffffff",
   19839 => x"ffffff",
   19840 => x"fffff5",
   19841 => x"c30c30",
   19842 => x"c30c30",
   19843 => x"c30c30",
   19844 => x"c30c30",
   19845 => x"c30c30",
   19846 => x"c30c30",
   19847 => x"c30c30",
   19848 => x"c30c30",
   19849 => x"c30c30",
   19850 => x"c30c30",
   19851 => x"c30c30",
   19852 => x"c30c30",
   19853 => x"c30c30",
   19854 => x"c30c30",
   19855 => x"c30c30",
   19856 => x"c30c30",
   19857 => x"c30c30",
   19858 => x"c219a7",
   19859 => x"df3cf3",
   19860 => x"cf3cf3",
   19861 => x"cf3cf3",
   19862 => x"cf3aae",
   19863 => x"ffffff",
   19864 => x"ffffff",
   19865 => x"ffffff",
   19866 => x"ffffff",
   19867 => x"ffffff",
   19868 => x"ffffff",
   19869 => x"ffffff",
   19870 => x"ffffff",
   19871 => x"ffffff",
   19872 => x"ffffff",
   19873 => x"ffffff",
   19874 => x"ffffff",
   19875 => x"ffffff",
   19876 => x"ffffff",
   19877 => x"ffffff",
   19878 => x"ffffff",
   19879 => x"ffffff",
   19880 => x"ffffff",
   19881 => x"ffffff",
   19882 => x"ffffff",
   19883 => x"ffffff",
   19884 => x"ffffff",
   19885 => x"ffffde",
   19886 => x"3cf3cf",
   19887 => x"3cf3cf",
   19888 => x"3cf3cf",
   19889 => x"3cf3ce",
   19890 => x"30c30c",
   19891 => x"30c30c",
   19892 => x"30c30c",
   19893 => x"30c30c",
   19894 => x"30c30c",
   19895 => x"30c30c",
   19896 => x"30c30c",
   19897 => x"30c30c",
   19898 => x"30c30c",
   19899 => x"30c30c",
   19900 => x"30c30c",
   19901 => x"30c30c",
   19902 => x"30c30c",
   19903 => x"30c30c",
   19904 => x"30c30c",
   19905 => x"30c30c",
   19906 => x"30c30c",
   19907 => x"30c32e",
   19908 => x"ffffff",
   19909 => x"ffffff",
   19910 => x"ffffff",
   19911 => x"ffffff",
   19912 => x"ffffff",
   19913 => x"ffffff",
   19914 => x"ffffff",
   19915 => x"ffffff",
   19916 => x"ffffff",
   19917 => x"ffffff",
   19918 => x"ffffff",
   19919 => x"ffffff",
   19920 => x"fffa95",
   19921 => x"abffff",
   19922 => x"ffffff",
   19923 => x"ffffff",
   19924 => x"ffffff",
   19925 => x"ffffff",
   19926 => x"ffffff",
   19927 => x"ffffff",
   19928 => x"ffffff",
   19929 => x"ffffff",
   19930 => x"ffffff",
   19931 => x"ffffff",
   19932 => x"ffffff",
   19933 => x"ffffff",
   19934 => x"ffffff",
   19935 => x"ffffff",
   19936 => x"ffffff",
   19937 => x"ffffff",
   19938 => x"ffffff",
   19939 => x"ffffff",
   19940 => x"ffffff",
   19941 => x"ffffff",
   19942 => x"ffffff",
   19943 => x"ffffff",
   19944 => x"ffffff",
   19945 => x"ffffff",
   19946 => x"ffffff",
   19947 => x"ffffff",
   19948 => x"ffffff",
   19949 => x"ffffff",
   19950 => x"ffffff",
   19951 => x"ffffff",
   19952 => x"ffffff",
   19953 => x"ffffff",
   19954 => x"ffffff",
   19955 => x"ffffff",
   19956 => x"ffffff",
   19957 => x"ffffff",
   19958 => x"ffffff",
   19959 => x"ffffff",
   19960 => x"ffffff",
   19961 => x"ffffff",
   19962 => x"ffffff",
   19963 => x"ffffff",
   19964 => x"ffffff",
   19965 => x"ffffff",
   19966 => x"ffffff",
   19967 => x"ffffff",
   19968 => x"ffffff",
   19969 => x"ffffff",
   19970 => x"ffffff",
   19971 => x"ffffff",
   19972 => x"ffffff",
   19973 => x"ffffff",
   19974 => x"ffffff",
   19975 => x"ffffff",
   19976 => x"ffffff",
   19977 => x"ffffff",
   19978 => x"ffffff",
   19979 => x"ffffff",
   19980 => x"ffffff",
   19981 => x"ffffff",
   19982 => x"ffffff",
   19983 => x"ffffff",
   19984 => x"ffffff",
   19985 => x"ffffff",
   19986 => x"ffffff",
   19987 => x"ffffff",
   19988 => x"ffffff",
   19989 => x"ffffff",
   19990 => x"ffffff",
   19991 => x"ffffff",
   19992 => x"ffffff",
   19993 => x"ffffff",
   19994 => x"ffffff",
   19995 => x"ffffff",
   19996 => x"ffffff",
   19997 => x"ffffff",
   19998 => x"ffffff",
   19999 => x"ffffff",
   20000 => x"fffffa",
   20001 => x"c30c30",
   20002 => x"c30c30",
   20003 => x"c30c30",
   20004 => x"c30c30",
   20005 => x"c30c30",
   20006 => x"c30c30",
   20007 => x"c30c30",
   20008 => x"c30c30",
   20009 => x"c30c30",
   20010 => x"c30c30",
   20011 => x"c30c30",
   20012 => x"c30c30",
   20013 => x"c30c30",
   20014 => x"c30c30",
   20015 => x"c30c30",
   20016 => x"c30c30",
   20017 => x"c30c30",
   20018 => x"8669f7",
   20019 => x"cf3cf3",
   20020 => x"cf3cf3",
   20021 => x"cf3cf3",
   20022 => x"cf39ae",
   20023 => x"ffffff",
   20024 => x"ffffff",
   20025 => x"ffffff",
   20026 => x"ffffff",
   20027 => x"ffffff",
   20028 => x"ffffff",
   20029 => x"ffffff",
   20030 => x"ffffff",
   20031 => x"ffffff",
   20032 => x"ffffff",
   20033 => x"ffffff",
   20034 => x"ffffff",
   20035 => x"ffffff",
   20036 => x"ffffff",
   20037 => x"ffffff",
   20038 => x"ffffff",
   20039 => x"ffffff",
   20040 => x"ffffff",
   20041 => x"ffffff",
   20042 => x"ffffff",
   20043 => x"ffffff",
   20044 => x"ffffff",
   20045 => x"ffffdd",
   20046 => x"3cf3cf",
   20047 => x"3cf3cf",
   20048 => x"3cf3cf",
   20049 => x"3cf3cf",
   20050 => x"38c30c",
   20051 => x"30c30c",
   20052 => x"30c30c",
   20053 => x"30c30c",
   20054 => x"30c30c",
   20055 => x"30c30c",
   20056 => x"30c30c",
   20057 => x"30c30c",
   20058 => x"30c30c",
   20059 => x"30c30c",
   20060 => x"30c30c",
   20061 => x"30c30c",
   20062 => x"30c30c",
   20063 => x"30c30c",
   20064 => x"30c30c",
   20065 => x"30c30c",
   20066 => x"30c30c",
   20067 => x"30c77f",
   20068 => x"ffffff",
   20069 => x"ffffff",
   20070 => x"ffffff",
   20071 => x"ffffff",
   20072 => x"ffffff",
   20073 => x"ffffff",
   20074 => x"ffffff",
   20075 => x"ffffff",
   20076 => x"ffffff",
   20077 => x"ffffff",
   20078 => x"ffffff",
   20079 => x"ffffff",
   20080 => x"fea56a",
   20081 => x"ffffff",
   20082 => x"ffffff",
   20083 => x"ffffff",
   20084 => x"ffffff",
   20085 => x"ffffff",
   20086 => x"ffffff",
   20087 => x"ffffff",
   20088 => x"ffffff",
   20089 => x"ffffff",
   20090 => x"ffffff",
   20091 => x"ffffff",
   20092 => x"ffffff",
   20093 => x"ffffff",
   20094 => x"ffffff",
   20095 => x"ffffff",
   20096 => x"ffffff",
   20097 => x"ffffff",
   20098 => x"ffffff",
   20099 => x"ffffff",
   20100 => x"ffffff",
   20101 => x"ffffff",
   20102 => x"ffffff",
   20103 => x"ffffff",
   20104 => x"ffffff",
   20105 => x"ffffff",
   20106 => x"ffffff",
   20107 => x"ffffff",
   20108 => x"ffffff",
   20109 => x"ffffff",
   20110 => x"ffffff",
   20111 => x"ffffff",
   20112 => x"ffffff",
   20113 => x"ffffff",
   20114 => x"ffffff",
   20115 => x"ffffff",
   20116 => x"ffffff",
   20117 => x"ffffff",
   20118 => x"ffffff",
   20119 => x"ffffff",
   20120 => x"ffffff",
   20121 => x"ffffff",
   20122 => x"ffffff",
   20123 => x"ffffff",
   20124 => x"ffffff",
   20125 => x"ffffff",
   20126 => x"ffffff",
   20127 => x"ffffff",
   20128 => x"ffffff",
   20129 => x"ffffff",
   20130 => x"ffffff",
   20131 => x"ffffff",
   20132 => x"ffffff",
   20133 => x"ffffff",
   20134 => x"ffffff",
   20135 => x"ffffff",
   20136 => x"ffffff",
   20137 => x"ffffff",
   20138 => x"ffffff",
   20139 => x"ffffff",
   20140 => x"ffffff",
   20141 => x"ffffff",
   20142 => x"ffffff",
   20143 => x"ffffff",
   20144 => x"ffffff",
   20145 => x"ffffff",
   20146 => x"ffffff",
   20147 => x"ffffff",
   20148 => x"ffffff",
   20149 => x"ffffff",
   20150 => x"ffffff",
   20151 => x"ffffff",
   20152 => x"ffffff",
   20153 => x"ffffff",
   20154 => x"ffffff",
   20155 => x"ffffff",
   20156 => x"ffffff",
   20157 => x"ffffff",
   20158 => x"ffffff",
   20159 => x"ffffff",
   20160 => x"ffffff",
   20161 => x"c30c30",
   20162 => x"c30c30",
   20163 => x"c30c30",
   20164 => x"c30c30",
   20165 => x"c30c30",
   20166 => x"c30c30",
   20167 => x"c30c30",
   20168 => x"c30c30",
   20169 => x"c30c30",
   20170 => x"c30c30",
   20171 => x"c30c30",
   20172 => x"c30c30",
   20173 => x"c30c30",
   20174 => x"c30c30",
   20175 => x"c30c30",
   20176 => x"c30c30",
   20177 => x"c30c21",
   20178 => x"5a7cf3",
   20179 => x"cf3cf3",
   20180 => x"cf3cf3",
   20181 => x"cf3cf3",
   20182 => x"cf39ea",
   20183 => x"bbffff",
   20184 => x"ffffff",
   20185 => x"ffffff",
   20186 => x"ffffff",
   20187 => x"ffffff",
   20188 => x"ffffff",
   20189 => x"ffffff",
   20190 => x"ffffff",
   20191 => x"ffffff",
   20192 => x"ffffff",
   20193 => x"ffffff",
   20194 => x"ffffff",
   20195 => x"ffffff",
   20196 => x"ffffff",
   20197 => x"ffffff",
   20198 => x"ffffff",
   20199 => x"ffffff",
   20200 => x"ffffff",
   20201 => x"ffffff",
   20202 => x"ffffff",
   20203 => x"ffffff",
   20204 => x"ffffff",
   20205 => x"fffb8d",
   20206 => x"3cf3cf",
   20207 => x"3cf3cf",
   20208 => x"3cf3cf",
   20209 => x"3cf3cf",
   20210 => x"3ce30c",
   20211 => x"30c30c",
   20212 => x"30c30c",
   20213 => x"30c30c",
   20214 => x"30c30c",
   20215 => x"30c30c",
   20216 => x"30c30c",
   20217 => x"30c30c",
   20218 => x"30c30c",
   20219 => x"30c30c",
   20220 => x"30c30c",
   20221 => x"30c30c",
   20222 => x"30c30c",
   20223 => x"30c30c",
   20224 => x"30c30c",
   20225 => x"30c30c",
   20226 => x"30c30c",
   20227 => x"30c77f",
   20228 => x"ffffff",
   20229 => x"ffffff",
   20230 => x"ffffff",
   20231 => x"ffffff",
   20232 => x"ffffff",
   20233 => x"ffffff",
   20234 => x"ffffff",
   20235 => x"ffffff",
   20236 => x"ffffff",
   20237 => x"ffffff",
   20238 => x"ffffff",
   20239 => x"ffffff",
   20240 => x"a95abf",
   20241 => x"ffffff",
   20242 => x"ffffff",
   20243 => x"ffffff",
   20244 => x"ffffff",
   20245 => x"ffffff",
   20246 => x"ffffff",
   20247 => x"ffffff",
   20248 => x"ffffff",
   20249 => x"ffffff",
   20250 => x"ffffff",
   20251 => x"ffffff",
   20252 => x"ffffff",
   20253 => x"ffffff",
   20254 => x"ffffff",
   20255 => x"ffffff",
   20256 => x"ffffff",
   20257 => x"ffffff",
   20258 => x"ffffff",
   20259 => x"ffffff",
   20260 => x"ffffff",
   20261 => x"ffffff",
   20262 => x"ffffff",
   20263 => x"ffffff",
   20264 => x"ffffff",
   20265 => x"ffffff",
   20266 => x"ffffff",
   20267 => x"ffffff",
   20268 => x"ffffff",
   20269 => x"ffffff",
   20270 => x"ffffff",
   20271 => x"ffffff",
   20272 => x"ffffff",
   20273 => x"ffffff",
   20274 => x"ffffff",
   20275 => x"ffffff",
   20276 => x"ffffff",
   20277 => x"ffffff",
   20278 => x"ffffff",
   20279 => x"ffffff",
   20280 => x"ffffff",
   20281 => x"ffffff",
   20282 => x"ffffff",
   20283 => x"ffffff",
   20284 => x"ffffff",
   20285 => x"ffffff",
   20286 => x"ffffff",
   20287 => x"ffffff",
   20288 => x"ffffff",
   20289 => x"ffffff",
   20290 => x"ffffff",
   20291 => x"ffffff",
   20292 => x"ffffff",
   20293 => x"ffffff",
   20294 => x"ffffff",
   20295 => x"ffffff",
   20296 => x"ffffff",
   20297 => x"ffffff",
   20298 => x"ffffff",
   20299 => x"ffffff",
   20300 => x"ffffff",
   20301 => x"ffffff",
   20302 => x"ffffff",
   20303 => x"ffffff",
   20304 => x"ffffff",
   20305 => x"ffffff",
   20306 => x"ffffff",
   20307 => x"ffffff",
   20308 => x"ffffff",
   20309 => x"ffffff",
   20310 => x"ffffff",
   20311 => x"ffffff",
   20312 => x"ffffff",
   20313 => x"ffffff",
   20314 => x"ffffff",
   20315 => x"ffffff",
   20316 => x"ffffff",
   20317 => x"ffffff",
   20318 => x"ffffff",
   20319 => x"ffffff",
   20320 => x"ffffff",
   20321 => x"d70c30",
   20322 => x"c30c30",
   20323 => x"c30c30",
   20324 => x"c30c30",
   20325 => x"c30c30",
   20326 => x"c30c30",
   20327 => x"c30c30",
   20328 => x"c30c30",
   20329 => x"c30c30",
   20330 => x"c30c30",
   20331 => x"c30c30",
   20332 => x"c30c30",
   20333 => x"c30c30",
   20334 => x"c30c30",
   20335 => x"c30c30",
   20336 => x"c30c30",
   20337 => x"c30866",
   20338 => x"9f3cf3",
   20339 => x"cf3cf3",
   20340 => x"cf3cf3",
   20341 => x"cf3cf3",
   20342 => x"cf3cea",
   20343 => x"bbffff",
   20344 => x"ffffff",
   20345 => x"ffffff",
   20346 => x"ffffff",
   20347 => x"ffffff",
   20348 => x"ffffff",
   20349 => x"ffffff",
   20350 => x"ffffff",
   20351 => x"ffffff",
   20352 => x"ffffff",
   20353 => x"ffffff",
   20354 => x"ffffff",
   20355 => x"ffffff",
   20356 => x"ffffff",
   20357 => x"ffffff",
   20358 => x"ffffff",
   20359 => x"ffffff",
   20360 => x"ffffff",
   20361 => x"ffffff",
   20362 => x"ffffff",
   20363 => x"ffffff",
   20364 => x"ffffff",
   20365 => x"fffb8e",
   20366 => x"3cf3cf",
   20367 => x"3cf3cf",
   20368 => x"3cf3cf",
   20369 => x"3cf3cf",
   20370 => x"3cf38c",
   20371 => x"30c30c",
   20372 => x"30c30c",
   20373 => x"30c30c",
   20374 => x"30c30c",
   20375 => x"30c30c",
   20376 => x"30c30c",
   20377 => x"30c30c",
   20378 => x"30c30c",
   20379 => x"30c30c",
   20380 => x"30c30c",
   20381 => x"30c30c",
   20382 => x"30c30c",
   20383 => x"30c30c",
   20384 => x"30c30c",
   20385 => x"30c30c",
   20386 => x"30c30c",
   20387 => x"30cbbf",
   20388 => x"ffffff",
   20389 => x"ffffff",
   20390 => x"ffffff",
   20391 => x"ffffff",
   20392 => x"ffffff",
   20393 => x"ffffff",
   20394 => x"ffffff",
   20395 => x"ffffff",
   20396 => x"ffffff",
   20397 => x"ffffff",
   20398 => x"ffffff",
   20399 => x"ffffea",
   20400 => x"56afff",
   20401 => x"ffffff",
   20402 => x"ffffff",
   20403 => x"ffffff",
   20404 => x"ffffff",
   20405 => x"ffffff",
   20406 => x"ffffff",
   20407 => x"ffffff",
   20408 => x"ffffff",
   20409 => x"ffffff",
   20410 => x"ffffff",
   20411 => x"ffffff",
   20412 => x"ffffff",
   20413 => x"ffffff",
   20414 => x"ffffff",
   20415 => x"ffffff",
   20416 => x"ffffff",
   20417 => x"ffffff",
   20418 => x"ffffff",
   20419 => x"ffffff",
   20420 => x"ffffff",
   20421 => x"ffffff",
   20422 => x"ffffff",
   20423 => x"ffffff",
   20424 => x"ffffff",
   20425 => x"ffffff",
   20426 => x"ffffff",
   20427 => x"ffffff",
   20428 => x"ffffff",
   20429 => x"ffffff",
   20430 => x"ffffff",
   20431 => x"ffffff",
   20432 => x"ffffff",
   20433 => x"ffffff",
   20434 => x"ffffff",
   20435 => x"ffffff",
   20436 => x"ffffff",
   20437 => x"ffffff",
   20438 => x"ffffff",
   20439 => x"ffffff",
   20440 => x"ffffff",
   20441 => x"ffffff",
   20442 => x"ffffff",
   20443 => x"ffffff",
   20444 => x"ffffff",
   20445 => x"ffffff",
   20446 => x"ffffff",
   20447 => x"ffffff",
   20448 => x"ffffff",
   20449 => x"ffffff",
   20450 => x"ffffff",
   20451 => x"ffffff",
   20452 => x"ffffff",
   20453 => x"ffffff",
   20454 => x"ffffff",
   20455 => x"ffffff",
   20456 => x"ffffff",
   20457 => x"ffffff",
   20458 => x"ffffff",
   20459 => x"ffffff",
   20460 => x"ffffff",
   20461 => x"ffffff",
   20462 => x"ffffff",
   20463 => x"ffffff",
   20464 => x"ffffff",
   20465 => x"ffffff",
   20466 => x"ffffff",
   20467 => x"ffffff",
   20468 => x"ffffff",
   20469 => x"ffffff",
   20470 => x"ffffff",
   20471 => x"ffffff",
   20472 => x"ffffff",
   20473 => x"ffffff",
   20474 => x"ffffff",
   20475 => x"ffffff",
   20476 => x"ffffff",
   20477 => x"ffffff",
   20478 => x"ffffff",
   20479 => x"ffffff",
   20480 => x"ffffff",
   20481 => x"d70c30",
   20482 => x"c30c30",
   20483 => x"c30c30",
   20484 => x"c30c30",
   20485 => x"c30c30",
   20486 => x"c30c30",
   20487 => x"c30c30",
   20488 => x"c30c30",
   20489 => x"c30c30",
   20490 => x"c30c30",
   20491 => x"c30c30",
   20492 => x"c30c30",
   20493 => x"c30c30",
   20494 => x"c30c30",
   20495 => x"c30c30",
   20496 => x"c30c30",
   20497 => x"c219a7",
   20498 => x"cf3cf3",
   20499 => x"cf3cf3",
   20500 => x"cf3cf3",
   20501 => x"cf3cf3",
   20502 => x"cf3ce6",
   20503 => x"bbffff",
   20504 => x"ffffff",
   20505 => x"ffffff",
   20506 => x"ffffff",
   20507 => x"ffffff",
   20508 => x"ffffff",
   20509 => x"ffffff",
   20510 => x"ffffff",
   20511 => x"ffffff",
   20512 => x"ffffff",
   20513 => x"ffffff",
   20514 => x"ffffff",
   20515 => x"ffffff",
   20516 => x"ffffff",
   20517 => x"ffffff",
   20518 => x"ffffff",
   20519 => x"ffffff",
   20520 => x"ffffff",
   20521 => x"ffffff",
   20522 => x"ffffff",
   20523 => x"ffffff",
   20524 => x"ffffff",
   20525 => x"fff78f",
   20526 => x"3cf3cf",
   20527 => x"3cf3cf",
   20528 => x"3cf3cf",
   20529 => x"3cf3cf",
   20530 => x"3cf3ce",
   20531 => x"30c30c",
   20532 => x"30c30c",
   20533 => x"30c30c",
   20534 => x"30c30c",
   20535 => x"30c30c",
   20536 => x"30c30c",
   20537 => x"30c30c",
   20538 => x"30c30c",
   20539 => x"30c30c",
   20540 => x"30c30c",
   20541 => x"30c30c",
   20542 => x"30c30c",
   20543 => x"30c30c",
   20544 => x"30c30c",
   20545 => x"30c30c",
   20546 => x"30c30c",
   20547 => x"30cbbf",
   20548 => x"ffffff",
   20549 => x"ffffff",
   20550 => x"ffffff",
   20551 => x"ffffff",
   20552 => x"ffffff",
   20553 => x"ffffff",
   20554 => x"ffffff",
   20555 => x"ffffff",
   20556 => x"ffffff",
   20557 => x"ffffff",
   20558 => x"ffffff",
   20559 => x"fffa95",
   20560 => x"abffff",
   20561 => x"ffffff",
   20562 => x"ffffff",
   20563 => x"ffffff",
   20564 => x"ffffff",
   20565 => x"ffffff",
   20566 => x"ffffff",
   20567 => x"ffffff",
   20568 => x"ffffff",
   20569 => x"ffffff",
   20570 => x"ffffff",
   20571 => x"ffffff",
   20572 => x"ffffff",
   20573 => x"ffffff",
   20574 => x"ffffff",
   20575 => x"ffffff",
   20576 => x"ffffff",
   20577 => x"ffffff",
   20578 => x"ffffff",
   20579 => x"ffffff",
   20580 => x"ffffff",
   20581 => x"ffffff",
   20582 => x"ffffff",
   20583 => x"ffffff",
   20584 => x"ffffff",
   20585 => x"ffffff",
   20586 => x"ffffff",
   20587 => x"ffffff",
   20588 => x"ffffff",
   20589 => x"ffffff",
   20590 => x"ffffff",
   20591 => x"ffffff",
   20592 => x"ffffff",
   20593 => x"ffffff",
   20594 => x"ffffff",
   20595 => x"ffffff",
   20596 => x"ffffff",
   20597 => x"ffffff",
   20598 => x"ffffff",
   20599 => x"ffffff",
   20600 => x"ffffff",
   20601 => x"ffffff",
   20602 => x"ffffff",
   20603 => x"ffffff",
   20604 => x"ffffff",
   20605 => x"ffffff",
   20606 => x"ffffff",
   20607 => x"ffffff",
   20608 => x"ffffff",
   20609 => x"ffffff",
   20610 => x"ffffff",
   20611 => x"ffffff",
   20612 => x"ffffff",
   20613 => x"ffffff",
   20614 => x"ffffff",
   20615 => x"ffffff",
   20616 => x"ffffff",
   20617 => x"ffffff",
   20618 => x"ffffff",
   20619 => x"ffffff",
   20620 => x"ffffff",
   20621 => x"ffffff",
   20622 => x"ffffff",
   20623 => x"ffffff",
   20624 => x"ffffff",
   20625 => x"ffffff",
   20626 => x"ffffff",
   20627 => x"ffffff",
   20628 => x"ffffff",
   20629 => x"ffffff",
   20630 => x"ffffff",
   20631 => x"ffffff",
   20632 => x"ffffff",
   20633 => x"ffffff",
   20634 => x"ffffff",
   20635 => x"ffffff",
   20636 => x"ffffff",
   20637 => x"ffffff",
   20638 => x"ffffff",
   20639 => x"ffffff",
   20640 => x"ffffff",
   20641 => x"eb0c30",
   20642 => x"c30c30",
   20643 => x"c30c30",
   20644 => x"c30c30",
   20645 => x"c30c30",
   20646 => x"c30c30",
   20647 => x"c30c30",
   20648 => x"c30c30",
   20649 => x"c30c30",
   20650 => x"c30c30",
   20651 => x"c30c30",
   20652 => x"c30c30",
   20653 => x"c30c30",
   20654 => x"c30c30",
   20655 => x"c30c30",
   20656 => x"c30c30",
   20657 => x"c669f3",
   20658 => x"cf3cf3",
   20659 => x"cf3cf3",
   20660 => x"cf3cf3",
   20661 => x"cf3cf3",
   20662 => x"cf3ce6",
   20663 => x"abffff",
   20664 => x"ffffff",
   20665 => x"ffffff",
   20666 => x"ffffff",
   20667 => x"ffffff",
   20668 => x"ffffff",
   20669 => x"ffffff",
   20670 => x"ffffff",
   20671 => x"ffffff",
   20672 => x"ffffff",
   20673 => x"ffffff",
   20674 => x"ffffff",
   20675 => x"ffffff",
   20676 => x"ffffff",
   20677 => x"ffffff",
   20678 => x"ffffff",
   20679 => x"ffffff",
   20680 => x"ffffff",
   20681 => x"ffffff",
   20682 => x"ffffff",
   20683 => x"ffffff",
   20684 => x"ffffff",
   20685 => x"fff34f",
   20686 => x"3cf3cf",
   20687 => x"3cf3cf",
   20688 => x"3cf3cf",
   20689 => x"3cf3cf",
   20690 => x"3cf3cf",
   20691 => x"38c30c",
   20692 => x"30c30c",
   20693 => x"30c30c",
   20694 => x"30c30c",
   20695 => x"30c30c",
   20696 => x"30c30c",
   20697 => x"30c30c",
   20698 => x"30c30c",
   20699 => x"30c30c",
   20700 => x"30c30c",
   20701 => x"30c30c",
   20702 => x"30c30c",
   20703 => x"30c30c",
   20704 => x"30c30c",
   20705 => x"30c30c",
   20706 => x"30c30c",
   20707 => x"31dfff",
   20708 => x"ffffff",
   20709 => x"ffffff",
   20710 => x"ffffff",
   20711 => x"ffffff",
   20712 => x"ffffff",
   20713 => x"ffffff",
   20714 => x"ffffff",
   20715 => x"ffffff",
   20716 => x"ffffff",
   20717 => x"ffffff",
   20718 => x"ffffff",
   20719 => x"fea56a",
   20720 => x"ffffff",
   20721 => x"ffffff",
   20722 => x"ffffff",
   20723 => x"ffffff",
   20724 => x"ffffff",
   20725 => x"ffffff",
   20726 => x"ffffff",
   20727 => x"ffffff",
   20728 => x"ffffff",
   20729 => x"ffffff",
   20730 => x"ffffff",
   20731 => x"ffffff",
   20732 => x"ffffff",
   20733 => x"ffffff",
   20734 => x"ffffff",
   20735 => x"ffffff",
   20736 => x"ffffff",
   20737 => x"ffffff",
   20738 => x"ffffff",
   20739 => x"ffffff",
   20740 => x"ffffff",
   20741 => x"ffffff",
   20742 => x"ffffff",
   20743 => x"ffffff",
   20744 => x"ffffff",
   20745 => x"ffffff",
   20746 => x"ffffff",
   20747 => x"ffffff",
   20748 => x"ffffff",
   20749 => x"ffffff",
   20750 => x"ffffff",
   20751 => x"ffffff",
   20752 => x"ffffff",
   20753 => x"ffffff",
   20754 => x"ffffff",
   20755 => x"ffffff",
   20756 => x"ffffff",
   20757 => x"ffffff",
   20758 => x"ffffff",
   20759 => x"ffffff",
   20760 => x"ffffff",
   20761 => x"ffffff",
   20762 => x"ffffff",
   20763 => x"ffffff",
   20764 => x"ffffff",
   20765 => x"ffffff",
   20766 => x"ffffff",
   20767 => x"ffffff",
   20768 => x"ffffff",
   20769 => x"ffffff",
   20770 => x"ffffff",
   20771 => x"ffffff",
   20772 => x"ffffff",
   20773 => x"ffffff",
   20774 => x"ffffff",
   20775 => x"ffffff",
   20776 => x"ffffff",
   20777 => x"ffffff",
   20778 => x"ffffff",
   20779 => x"ffffff",
   20780 => x"ffffff",
   20781 => x"ffffff",
   20782 => x"ffffff",
   20783 => x"ffffff",
   20784 => x"ffffff",
   20785 => x"ffffff",
   20786 => x"ffffff",
   20787 => x"ffffff",
   20788 => x"ffffff",
   20789 => x"ffffff",
   20790 => x"ffffff",
   20791 => x"ffffff",
   20792 => x"ffffff",
   20793 => x"ffffff",
   20794 => x"ffffff",
   20795 => x"ffffff",
   20796 => x"ffffff",
   20797 => x"ffffff",
   20798 => x"ffffff",
   20799 => x"ffffff",
   20800 => x"ffffff",
   20801 => x"ff5c30",
   20802 => x"c30c30",
   20803 => x"c30c30",
   20804 => x"c30c30",
   20805 => x"c30c30",
   20806 => x"c30c30",
   20807 => x"c30c30",
   20808 => x"c30c30",
   20809 => x"c30c30",
   20810 => x"c30c30",
   20811 => x"c30c30",
   20812 => x"c30c30",
   20813 => x"c30c30",
   20814 => x"c30c30",
   20815 => x"c30c30",
   20816 => x"c30c30",
   20817 => x"9a7df3",
   20818 => x"cf3cf3",
   20819 => x"cf3cf3",
   20820 => x"cf3cf3",
   20821 => x"cf3cf3",
   20822 => x"cf3cf3",
   20823 => x"abefff",
   20824 => x"ffffff",
   20825 => x"ffffff",
   20826 => x"ffffff",
   20827 => x"ffffff",
   20828 => x"ffffff",
   20829 => x"ffffff",
   20830 => x"ffffff",
   20831 => x"ffffff",
   20832 => x"ffffff",
   20833 => x"ffffff",
   20834 => x"ffffff",
   20835 => x"ffffff",
   20836 => x"ffffff",
   20837 => x"ffffff",
   20838 => x"ffffff",
   20839 => x"ffffff",
   20840 => x"ffffff",
   20841 => x"ffffff",
   20842 => x"ffffff",
   20843 => x"ffffff",
   20844 => x"ffffff",
   20845 => x"fee38f",
   20846 => x"3cf3cf",
   20847 => x"3cf3cf",
   20848 => x"3cf3cf",
   20849 => x"3cf3cf",
   20850 => x"3cf3cf",
   20851 => x"3ce30c",
   20852 => x"30c30c",
   20853 => x"30c30c",
   20854 => x"30c30c",
   20855 => x"30c30c",
   20856 => x"30c30c",
   20857 => x"30c30c",
   20858 => x"30c30c",
   20859 => x"30c30c",
   20860 => x"30c30c",
   20861 => x"30c30c",
   20862 => x"30c30c",
   20863 => x"30c30c",
   20864 => x"30c30c",
   20865 => x"30c30c",
   20866 => x"30c30c",
   20867 => x"31dfff",
   20868 => x"ffffff",
   20869 => x"ffffff",
   20870 => x"ffffff",
   20871 => x"ffffff",
   20872 => x"ffffff",
   20873 => x"ffffff",
   20874 => x"ffffff",
   20875 => x"ffffff",
   20876 => x"ffffff",
   20877 => x"ffffff",
   20878 => x"ffffff",
   20879 => x"a95abf",
   20880 => x"ffffff",
   20881 => x"fffeb5",
   20882 => x"c30c30",
   20883 => x"c30c30",
   20884 => x"c30c30",
   20885 => x"c30c30",
   20886 => x"c30c30",
   20887 => x"c30c30",
   20888 => x"c30c30",
   20889 => x"c30c30",
   20890 => x"c30c30",
   20891 => x"c30c30",
   20892 => x"c30c30",
   20893 => x"c30c30",
   20894 => x"c30c30",
   20895 => x"820820",
   20896 => x"820820",
   20897 => x"820820",
   20898 => x"820820",
   20899 => x"820820",
   20900 => x"820820",
   20901 => x"820820",
   20902 => x"820820",
   20903 => x"820820",
   20904 => x"820820",
   20905 => x"820820",
   20906 => x"820820",
   20907 => x"820820",
   20908 => x"820820",
   20909 => x"820820",
   20910 => x"820820",
   20911 => x"820820",
   20912 => x"820820",
   20913 => x"820820",
   20914 => x"820820",
   20915 => x"820820",
   20916 => x"820820",
   20917 => x"820820",
   20918 => x"820820",
   20919 => x"820820",
   20920 => x"820820",
   20921 => x"820410",
   20922 => x"410410",
   20923 => x"410410",
   20924 => x"410410",
   20925 => x"410410",
   20926 => x"410410",
   20927 => x"410410",
   20928 => x"410410",
   20929 => x"410410",
   20930 => x"410410",
   20931 => x"410410",
   20932 => x"410410",
   20933 => x"410410",
   20934 => x"410410",
   20935 => x"410410",
   20936 => x"410410",
   20937 => x"410410",
   20938 => x"410410",
   20939 => x"410410",
   20940 => x"410410",
   20941 => x"410410",
   20942 => x"410410",
   20943 => x"410410",
   20944 => x"410410",
   20945 => x"410410",
   20946 => x"410410",
   20947 => x"410410",
   20948 => x"400000",
   20949 => x"000abf",
   20950 => x"ffffff",
   20951 => x"ffffff",
   20952 => x"ffffff",
   20953 => x"ffffff",
   20954 => x"ffffff",
   20955 => x"ffffff",
   20956 => x"ffffff",
   20957 => x"ffffff",
   20958 => x"ffffff",
   20959 => x"ffffff",
   20960 => x"ffffff",
   20961 => x"ff5c30",
   20962 => x"c30c30",
   20963 => x"c30c30",
   20964 => x"c30c30",
   20965 => x"c30c30",
   20966 => x"c30c30",
   20967 => x"c30c30",
   20968 => x"c30c30",
   20969 => x"c30c30",
   20970 => x"c30c30",
   20971 => x"c30c30",
   20972 => x"c30c30",
   20973 => x"c30c30",
   20974 => x"c30c30",
   20975 => x"c30c30",
   20976 => x"c30c26",
   20977 => x"9f7cf3",
   20978 => x"cf3cf3",
   20979 => x"cf3cf3",
   20980 => x"cf3cf3",
   20981 => x"cf3cf3",
   20982 => x"cf3cf3",
   20983 => x"aaefff",
   20984 => x"ffffff",
   20985 => x"ffffff",
   20986 => x"ffffff",
   20987 => x"ffffff",
   20988 => x"ffffff",
   20989 => x"ffffff",
   20990 => x"ffffff",
   20991 => x"ffffff",
   20992 => x"ffffff",
   20993 => x"ffffff",
   20994 => x"ffffff",
   20995 => x"ffffff",
   20996 => x"ffffff",
   20997 => x"ffffff",
   20998 => x"ffffff",
   20999 => x"ffffff",
   21000 => x"ffffff",
   21001 => x"ffffff",
   21002 => x"ffffff",
   21003 => x"ffffff",
   21004 => x"ffffff",
   21005 => x"fee38f",
   21006 => x"3cf3cf",
   21007 => x"3cf3cf",
   21008 => x"3cf3cf",
   21009 => x"3cf3cf",
   21010 => x"3cf3cf",
   21011 => x"3cf38c",
   21012 => x"30c30c",
   21013 => x"30c30c",
   21014 => x"30c30c",
   21015 => x"30c30c",
   21016 => x"30c30c",
   21017 => x"30c30c",
   21018 => x"30c30c",
   21019 => x"30c30c",
   21020 => x"30c30c",
   21021 => x"30c30c",
   21022 => x"30c30c",
   21023 => x"30c30c",
   21024 => x"30c30c",
   21025 => x"30c30c",
   21026 => x"30c30c",
   21027 => x"32efff",
   21028 => x"ffffff",
   21029 => x"ffffff",
   21030 => x"ffffff",
   21031 => x"ffffff",
   21032 => x"ffffff",
   21033 => x"ffffff",
   21034 => x"ffffff",
   21035 => x"ffffff",
   21036 => x"ffffff",
   21037 => x"ffffff",
   21038 => x"ffffea",
   21039 => x"56afff",
   21040 => x"ffffff",
   21041 => x"fffeb0",
   21042 => x"c30c30",
   21043 => x"c30c30",
   21044 => x"c30c30",
   21045 => x"c30c30",
   21046 => x"c30c30",
   21047 => x"c30c30",
   21048 => x"c30c30",
   21049 => x"c30c30",
   21050 => x"c30c30",
   21051 => x"c30c30",
   21052 => x"c30c30",
   21053 => x"820820",
   21054 => x"820820",
   21055 => x"820820",
   21056 => x"820820",
   21057 => x"820820",
   21058 => x"820820",
   21059 => x"820820",
   21060 => x"820820",
   21061 => x"820820",
   21062 => x"820820",
   21063 => x"820820",
   21064 => x"820820",
   21065 => x"820820",
   21066 => x"820820",
   21067 => x"820820",
   21068 => x"820820",
   21069 => x"820820",
   21070 => x"820820",
   21071 => x"820820",
   21072 => x"820820",
   21073 => x"820820",
   21074 => x"820820",
   21075 => x"820810",
   21076 => x"410410",
   21077 => x"410410",
   21078 => x"410410",
   21079 => x"410410",
   21080 => x"410410",
   21081 => x"410410",
   21082 => x"410410",
   21083 => x"410410",
   21084 => x"410410",
   21085 => x"410410",
   21086 => x"410410",
   21087 => x"410410",
   21088 => x"410410",
   21089 => x"410410",
   21090 => x"410410",
   21091 => x"410410",
   21092 => x"410410",
   21093 => x"410410",
   21094 => x"410410",
   21095 => x"410410",
   21096 => x"410410",
   21097 => x"410410",
   21098 => x"410400",
   21099 => x"000000",
   21100 => x"000000",
   21101 => x"000000",
   21102 => x"000000",
   21103 => x"000000",
   21104 => x"000000",
   21105 => x"000000",
   21106 => x"000000",
   21107 => x"000000",
   21108 => x"000000",
   21109 => x"00057f",
   21110 => x"ffffff",
   21111 => x"ffffff",
   21112 => x"ffffff",
   21113 => x"ffffff",
   21114 => x"ffffff",
   21115 => x"ffffff",
   21116 => x"ffffff",
   21117 => x"ffffff",
   21118 => x"ffffff",
   21119 => x"ffffff",
   21120 => x"ffffff",
   21121 => x"ffac30",
   21122 => x"c30c30",
   21123 => x"c30c30",
   21124 => x"c30c30",
   21125 => x"c30c30",
   21126 => x"c30c30",
   21127 => x"c30c30",
   21128 => x"c30c30",
   21129 => x"c30c30",
   21130 => x"c30c30",
   21131 => x"c30c30",
   21132 => x"c30c30",
   21133 => x"c30c30",
   21134 => x"c30c30",
   21135 => x"c30c30",
   21136 => x"c308a7",
   21137 => x"df3cf3",
   21138 => x"cf3cf3",
   21139 => x"cf3cf3",
   21140 => x"cf3cf3",
   21141 => x"cf3cf3",
   21142 => x"cf3cf3",
   21143 => x"9aefff",
   21144 => x"ffffff",
   21145 => x"ffffff",
   21146 => x"ffffff",
   21147 => x"ffffff",
   21148 => x"ffffff",
   21149 => x"ffffff",
   21150 => x"ffffff",
   21151 => x"ffffff",
   21152 => x"ffffff",
   21153 => x"ffffff",
   21154 => x"ffffff",
   21155 => x"ffffff",
   21156 => x"ffffff",
   21157 => x"ffffff",
   21158 => x"ffffff",
   21159 => x"ffffff",
   21160 => x"ffffff",
   21161 => x"ffffff",
   21162 => x"ffffff",
   21163 => x"ffffff",
   21164 => x"ffffff",
   21165 => x"fde3cf",
   21166 => x"3cf3cf",
   21167 => x"3cf3cf",
   21168 => x"3cf3cf",
   21169 => x"3cf3cf",
   21170 => x"3cf3cf",
   21171 => x"3cf3cd",
   21172 => x"30c30c",
   21173 => x"30c30c",
   21174 => x"30c30c",
   21175 => x"30c30c",
   21176 => x"30c30c",
   21177 => x"30c30c",
   21178 => x"30c30c",
   21179 => x"30c30c",
   21180 => x"30c30c",
   21181 => x"30c30c",
   21182 => x"30c30c",
   21183 => x"30c30c",
   21184 => x"30c30c",
   21185 => x"30c30c",
   21186 => x"30c30c",
   21187 => x"33ffff",
   21188 => x"ffffff",
   21189 => x"ffffff",
   21190 => x"ffffff",
   21191 => x"ffffff",
   21192 => x"ffffff",
   21193 => x"ffffff",
   21194 => x"ffffff",
   21195 => x"ffffff",
   21196 => x"ffffff",
   21197 => x"ffffff",
   21198 => x"fffa95",
   21199 => x"abffff",
   21200 => x"ffffff",
   21201 => x"fffeb0",
   21202 => x"c30c30",
   21203 => x"c30c30",
   21204 => x"c30c30",
   21205 => x"c30c30",
   21206 => x"c30c30",
   21207 => x"c30c30",
   21208 => x"c30c30",
   21209 => x"c30c30",
   21210 => x"c30c30",
   21211 => x"c30c30",
   21212 => x"c30c30",
   21213 => x"820820",
   21214 => x"820820",
   21215 => x"820820",
   21216 => x"820820",
   21217 => x"820820",
   21218 => x"820820",
   21219 => x"820820",
   21220 => x"820820",
   21221 => x"820820",
   21222 => x"820820",
   21223 => x"820820",
   21224 => x"820820",
   21225 => x"820820",
   21226 => x"820820",
   21227 => x"820820",
   21228 => x"820820",
   21229 => x"820820",
   21230 => x"820820",
   21231 => x"820820",
   21232 => x"820820",
   21233 => x"820820",
   21234 => x"820820",
   21235 => x"820410",
   21236 => x"410410",
   21237 => x"410410",
   21238 => x"410410",
   21239 => x"410410",
   21240 => x"410410",
   21241 => x"410410",
   21242 => x"410410",
   21243 => x"410410",
   21244 => x"410410",
   21245 => x"410410",
   21246 => x"410410",
   21247 => x"410410",
   21248 => x"410410",
   21249 => x"410410",
   21250 => x"410410",
   21251 => x"410410",
   21252 => x"410410",
   21253 => x"410410",
   21254 => x"410410",
   21255 => x"410410",
   21256 => x"410410",
   21257 => x"410410",
   21258 => x"410000",
   21259 => x"000000",
   21260 => x"000000",
   21261 => x"000000",
   21262 => x"000000",
   21263 => x"000000",
   21264 => x"000000",
   21265 => x"000000",
   21266 => x"000000",
   21267 => x"000000",
   21268 => x"000000",
   21269 => x"00057f",
   21270 => x"ffffff",
   21271 => x"ffffff",
   21272 => x"ffffff",
   21273 => x"ffffff",
   21274 => x"ffffff",
   21275 => x"ffffff",
   21276 => x"ffffff",
   21277 => x"ffffff",
   21278 => x"ffffff",
   21279 => x"ffffff",
   21280 => x"ffffff",
   21281 => x"ffac30",
   21282 => x"c30c30",
   21283 => x"c30c30",
   21284 => x"c30c30",
   21285 => x"c30c30",
   21286 => x"c30c30",
   21287 => x"c30c30",
   21288 => x"c30c30",
   21289 => x"c30c30",
   21290 => x"c30c30",
   21291 => x"c30c30",
   21292 => x"c30c30",
   21293 => x"c30c30",
   21294 => x"c30c30",
   21295 => x"c30c30",
   21296 => x"c219f7",
   21297 => x"cf3cf3",
   21298 => x"cf3cf3",
   21299 => x"cf3cf3",
   21300 => x"cf3cf3",
   21301 => x"cf3cf3",
   21302 => x"cf3cf3",
   21303 => x"9ebfff",
   21304 => x"ffffff",
   21305 => x"ffffff",
   21306 => x"ffffff",
   21307 => x"ffffff",
   21308 => x"ffffff",
   21309 => x"ffffff",
   21310 => x"ffffff",
   21311 => x"ffffff",
   21312 => x"ffffff",
   21313 => x"ffffff",
   21314 => x"ffffff",
   21315 => x"ffffff",
   21316 => x"ffffff",
   21317 => x"ffffff",
   21318 => x"ffffff",
   21319 => x"ffffff",
   21320 => x"ffffff",
   21321 => x"ffffff",
   21322 => x"ffffff",
   21323 => x"ffffff",
   21324 => x"ffffff",
   21325 => x"bce3cf",
   21326 => x"3cf3cf",
   21327 => x"3cf3cf",
   21328 => x"3cf3cf",
   21329 => x"3cf3cf",
   21330 => x"3cf3cf",
   21331 => x"3cf3ce",
   21332 => x"34c30c",
   21333 => x"30c30c",
   21334 => x"30c30c",
   21335 => x"30c30c",
   21336 => x"30c30c",
   21337 => x"30c30c",
   21338 => x"30c30c",
   21339 => x"30c30c",
   21340 => x"30c30c",
   21341 => x"30c30c",
   21342 => x"30c30c",
   21343 => x"30c30c",
   21344 => x"30c30c",
   21345 => x"30c30c",
   21346 => x"30c30c",
   21347 => x"77ffff",
   21348 => x"ffffff",
   21349 => x"ffffff",
   21350 => x"ffffff",
   21351 => x"ffffff",
   21352 => x"ffffff",
   21353 => x"ffffff",
   21354 => x"ffffff",
   21355 => x"ffffff",
   21356 => x"ffffff",
   21357 => x"ffffff",
   21358 => x"fea56a",
   21359 => x"ffffff",
   21360 => x"ffffff",
   21361 => x"fffeb0",
   21362 => x"c30c30",
   21363 => x"c30c30",
   21364 => x"c30c30",
   21365 => x"c30c30",
   21366 => x"c30c30",
   21367 => x"c30c30",
   21368 => x"c30c30",
   21369 => x"c30c30",
   21370 => x"c30c30",
   21371 => x"c30c30",
   21372 => x"c30c30",
   21373 => x"820820",
   21374 => x"820820",
   21375 => x"820820",
   21376 => x"820820",
   21377 => x"820820",
   21378 => x"820820",
   21379 => x"820820",
   21380 => x"820820",
   21381 => x"820820",
   21382 => x"820820",
   21383 => x"820820",
   21384 => x"820820",
   21385 => x"820820",
   21386 => x"820820",
   21387 => x"820820",
   21388 => x"820820",
   21389 => x"820820",
   21390 => x"820820",
   21391 => x"820820",
   21392 => x"820820",
   21393 => x"820820",
   21394 => x"820820",
   21395 => x"820410",
   21396 => x"410410",
   21397 => x"410410",
   21398 => x"410410",
   21399 => x"410410",
   21400 => x"410410",
   21401 => x"410410",
   21402 => x"410410",
   21403 => x"410410",
   21404 => x"410410",
   21405 => x"410410",
   21406 => x"410410",
   21407 => x"410410",
   21408 => x"410410",
   21409 => x"410410",
   21410 => x"410410",
   21411 => x"410410",
   21412 => x"410410",
   21413 => x"410410",
   21414 => x"410410",
   21415 => x"410410",
   21416 => x"410410",
   21417 => x"410410",
   21418 => x"410000",
   21419 => x"000000",
   21420 => x"000000",
   21421 => x"000000",
   21422 => x"000000",
   21423 => x"000000",
   21424 => x"000000",
   21425 => x"000000",
   21426 => x"000000",
   21427 => x"000000",
   21428 => x"000000",
   21429 => x"00057f",
   21430 => x"ffffff",
   21431 => x"ffffff",
   21432 => x"ffffff",
   21433 => x"ffffff",
   21434 => x"ffffff",
   21435 => x"ffffff",
   21436 => x"ffffff",
   21437 => x"ffffff",
   21438 => x"ffffff",
   21439 => x"ffffff",
   21440 => x"ffffff",
   21441 => x"fffd70",
   21442 => x"c30c30",
   21443 => x"c30c30",
   21444 => x"c30c30",
   21445 => x"c30c30",
   21446 => x"c30c30",
   21447 => x"c30c30",
   21448 => x"c30c30",
   21449 => x"c30c30",
   21450 => x"c30c30",
   21451 => x"c30c30",
   21452 => x"c30c30",
   21453 => x"c30c30",
   21454 => x"c30c30",
   21455 => x"c30c30",
   21456 => x"866df3",
   21457 => x"cf3cf3",
   21458 => x"cf3cf3",
   21459 => x"cf3cf3",
   21460 => x"cf3cf3",
   21461 => x"cf3cf3",
   21462 => x"cf3cf3",
   21463 => x"deabbf",
   21464 => x"ffffff",
   21465 => x"ffffff",
   21466 => x"ffffff",
   21467 => x"ffffff",
   21468 => x"ffffff",
   21469 => x"ffffff",
   21470 => x"ffffff",
   21471 => x"ffffff",
   21472 => x"ffffff",
   21473 => x"ffffff",
   21474 => x"ffffff",
   21475 => x"ffffff",
   21476 => x"ffffff",
   21477 => x"ffffff",
   21478 => x"ffffff",
   21479 => x"ffffff",
   21480 => x"ffffff",
   21481 => x"ffffff",
   21482 => x"ffffff",
   21483 => x"ffffff",
   21484 => x"ffffff",
   21485 => x"b8e3cf",
   21486 => x"3cf3cf",
   21487 => x"3cf3cf",
   21488 => x"3cf3cf",
   21489 => x"3cf3cf",
   21490 => x"3cf3cf",
   21491 => x"3cf3cf",
   21492 => x"38d30c",
   21493 => x"30c30c",
   21494 => x"30c30c",
   21495 => x"30c30c",
   21496 => x"30c30c",
   21497 => x"30c30c",
   21498 => x"30c30c",
   21499 => x"30c30c",
   21500 => x"30c30c",
   21501 => x"30c30c",
   21502 => x"30c30c",
   21503 => x"30c30c",
   21504 => x"30c30c",
   21505 => x"30c30c",
   21506 => x"30c30c",
   21507 => x"bbffff",
   21508 => x"ffffff",
   21509 => x"ffffff",
   21510 => x"ffffff",
   21511 => x"ffffff",
   21512 => x"ffffff",
   21513 => x"ffffff",
   21514 => x"ffffff",
   21515 => x"ffffff",
   21516 => x"ffffff",
   21517 => x"ffffff",
   21518 => x"a95abf",
   21519 => x"ffffff",
   21520 => x"ffffff",
   21521 => x"fffeb0",
   21522 => x"c30c30",
   21523 => x"c30c30",
   21524 => x"c30c30",
   21525 => x"c30c30",
   21526 => x"c30c30",
   21527 => x"c30c30",
   21528 => x"c30c30",
   21529 => x"c30c30",
   21530 => x"c30c30",
   21531 => x"c30c30",
   21532 => x"c30c30",
   21533 => x"820820",
   21534 => x"820820",
   21535 => x"820820",
   21536 => x"820820",
   21537 => x"820820",
   21538 => x"820820",
   21539 => x"820820",
   21540 => x"820820",
   21541 => x"820820",
   21542 => x"820820",
   21543 => x"820820",
   21544 => x"820820",
   21545 => x"820820",
   21546 => x"820820",
   21547 => x"820820",
   21548 => x"820820",
   21549 => x"820820",
   21550 => x"820820",
   21551 => x"820820",
   21552 => x"820820",
   21553 => x"820820",
   21554 => x"820820",
   21555 => x"820410",
   21556 => x"410410",
   21557 => x"410410",
   21558 => x"410410",
   21559 => x"410410",
   21560 => x"410410",
   21561 => x"410410",
   21562 => x"410410",
   21563 => x"410410",
   21564 => x"410410",
   21565 => x"410410",
   21566 => x"410410",
   21567 => x"410410",
   21568 => x"410410",
   21569 => x"410410",
   21570 => x"410410",
   21571 => x"410410",
   21572 => x"410410",
   21573 => x"410410",
   21574 => x"410410",
   21575 => x"410410",
   21576 => x"410410",
   21577 => x"410410",
   21578 => x"410000",
   21579 => x"000000",
   21580 => x"000000",
   21581 => x"000000",
   21582 => x"000000",
   21583 => x"000000",
   21584 => x"000000",
   21585 => x"000000",
   21586 => x"000000",
   21587 => x"000000",
   21588 => x"000000",
   21589 => x"00057f",
   21590 => x"ffffff",
   21591 => x"ffffff",
   21592 => x"ffffff",
   21593 => x"ffffff",
   21594 => x"ffffff",
   21595 => x"ffffff",
   21596 => x"ffffff",
   21597 => x"ffffff",
   21598 => x"ffffff",
   21599 => x"ffffff",
   21600 => x"ffffff",
   21601 => x"fffeb0",
   21602 => x"c30c30",
   21603 => x"c30c30",
   21604 => x"c30c30",
   21605 => x"c30c30",
   21606 => x"c30c30",
   21607 => x"c30c30",
   21608 => x"c30c30",
   21609 => x"c30c30",
   21610 => x"c30c30",
   21611 => x"c30c30",
   21612 => x"c30c30",
   21613 => x"c30c30",
   21614 => x"c30c30",
   21615 => x"c30c21",
   21616 => x"9a7cf3",
   21617 => x"cf3cf3",
   21618 => x"cf3cf3",
   21619 => x"cf3cf3",
   21620 => x"cf3cf3",
   21621 => x"cf3cf3",
   21622 => x"cf3cf3",
   21623 => x"ce6bbf",
   21624 => x"ffffff",
   21625 => x"ffffff",
   21626 => x"ffffff",
   21627 => x"ffffff",
   21628 => x"ffffff",
   21629 => x"ffffff",
   21630 => x"ffffff",
   21631 => x"ffffff",
   21632 => x"ffffff",
   21633 => x"ffffff",
   21634 => x"ffffff",
   21635 => x"ffffff",
   21636 => x"ffffff",
   21637 => x"ffffff",
   21638 => x"ffffff",
   21639 => x"ffffff",
   21640 => x"ffffff",
   21641 => x"ffffff",
   21642 => x"ffffff",
   21643 => x"ffffff",
   21644 => x"ffffff",
   21645 => x"78f3cf",
   21646 => x"3cf3cf",
   21647 => x"3cf3cf",
   21648 => x"3cf3cf",
   21649 => x"3cf3cf",
   21650 => x"3cf3cf",
   21651 => x"3cf3cf",
   21652 => x"3ce30c",
   21653 => x"30c30c",
   21654 => x"30c30c",
   21655 => x"30c30c",
   21656 => x"30c30c",
   21657 => x"30c30c",
   21658 => x"30c30c",
   21659 => x"30c30c",
   21660 => x"30c30c",
   21661 => x"30c30c",
   21662 => x"30c30c",
   21663 => x"30c30c",
   21664 => x"30c30c",
   21665 => x"30c30c",
   21666 => x"30c30c",
   21667 => x"ffffff",
   21668 => x"ffffff",
   21669 => x"ffffff",
   21670 => x"ffffff",
   21671 => x"ffffff",
   21672 => x"ffffff",
   21673 => x"ffffff",
   21674 => x"ffffff",
   21675 => x"ffffff",
   21676 => x"ffffff",
   21677 => x"ffffea",
   21678 => x"56afff",
   21679 => x"ffffff",
   21680 => x"ffffff",
   21681 => x"fffeb0",
   21682 => x"c30c30",
   21683 => x"c30c30",
   21684 => x"c30c30",
   21685 => x"c30c30",
   21686 => x"c30c30",
   21687 => x"c30c30",
   21688 => x"c30c30",
   21689 => x"c30c30",
   21690 => x"c30c30",
   21691 => x"c30c30",
   21692 => x"c30c30",
   21693 => x"820820",
   21694 => x"820820",
   21695 => x"820820",
   21696 => x"820820",
   21697 => x"820820",
   21698 => x"820820",
   21699 => x"820820",
   21700 => x"820820",
   21701 => x"820820",
   21702 => x"820820",
   21703 => x"820820",
   21704 => x"820820",
   21705 => x"820820",
   21706 => x"820820",
   21707 => x"820820",
   21708 => x"820820",
   21709 => x"820820",
   21710 => x"820820",
   21711 => x"820820",
   21712 => x"820820",
   21713 => x"820820",
   21714 => x"820820",
   21715 => x"820410",
   21716 => x"410410",
   21717 => x"410410",
   21718 => x"410410",
   21719 => x"410410",
   21720 => x"410410",
   21721 => x"410410",
   21722 => x"410410",
   21723 => x"410410",
   21724 => x"410410",
   21725 => x"410410",
   21726 => x"410410",
   21727 => x"410410",
   21728 => x"410410",
   21729 => x"410410",
   21730 => x"410410",
   21731 => x"410410",
   21732 => x"410410",
   21733 => x"410410",
   21734 => x"410410",
   21735 => x"410410",
   21736 => x"410410",
   21737 => x"410410",
   21738 => x"410000",
   21739 => x"000000",
   21740 => x"000000",
   21741 => x"000000",
   21742 => x"000000",
   21743 => x"000000",
   21744 => x"000000",
   21745 => x"000000",
   21746 => x"000000",
   21747 => x"000000",
   21748 => x"000000",
   21749 => x"00057f",
   21750 => x"ffffff",
   21751 => x"ffffff",
   21752 => x"ffffff",
   21753 => x"ffffff",
   21754 => x"ffffff",
   21755 => x"ffffff",
   21756 => x"ffffff",
   21757 => x"ffffff",
   21758 => x"ffffff",
   21759 => x"ffffff",
   21760 => x"ffffff",
   21761 => x"fffff5",
   21762 => x"c30c30",
   21763 => x"c30c30",
   21764 => x"c30c30",
   21765 => x"c30c30",
   21766 => x"c30c30",
   21767 => x"c30c30",
   21768 => x"c30c30",
   21769 => x"c30c30",
   21770 => x"c30c30",
   21771 => x"c30c30",
   21772 => x"c30c30",
   21773 => x"c30c30",
   21774 => x"c30c30",
   21775 => x"c30c22",
   21776 => x"9f3cf3",
   21777 => x"cf3cf3",
   21778 => x"cf3cf3",
   21779 => x"cf3cf3",
   21780 => x"cf3cf3",
   21781 => x"cf3cf3",
   21782 => x"cf3cf3",
   21783 => x"ce7abf",
   21784 => x"ffffff",
   21785 => x"ffffff",
   21786 => x"ffffff",
   21787 => x"ffffff",
   21788 => x"ffffff",
   21789 => x"ffffff",
   21790 => x"ffffff",
   21791 => x"ffffff",
   21792 => x"ffffff",
   21793 => x"ffffff",
   21794 => x"ffffff",
   21795 => x"ffffff",
   21796 => x"ffffff",
   21797 => x"ffffff",
   21798 => x"ffffff",
   21799 => x"ffffff",
   21800 => x"ffffff",
   21801 => x"ffffff",
   21802 => x"ffffff",
   21803 => x"ffffff",
   21804 => x"ffffee",
   21805 => x"34f3cf",
   21806 => x"3cf3cf",
   21807 => x"3cf3cf",
   21808 => x"3cf3cf",
   21809 => x"3cf3cf",
   21810 => x"3cf3cf",
   21811 => x"3cf3cf",
   21812 => x"3cf38c",
   21813 => x"30c30c",
   21814 => x"30c30c",
   21815 => x"30c30c",
   21816 => x"30c30c",
   21817 => x"30c30c",
   21818 => x"30c30c",
   21819 => x"30c30c",
   21820 => x"30c30c",
   21821 => x"30c30c",
   21822 => x"30c30c",
   21823 => x"30c30c",
   21824 => x"30c30c",
   21825 => x"30c30c",
   21826 => x"30c31d",
   21827 => x"ffffff",
   21828 => x"ffffff",
   21829 => x"ffffff",
   21830 => x"ffffff",
   21831 => x"ffffff",
   21832 => x"ffffff",
   21833 => x"ffffff",
   21834 => x"ffffff",
   21835 => x"ffffff",
   21836 => x"ffffff",
   21837 => x"fffa95",
   21838 => x"abffff",
   21839 => x"ffffff",
   21840 => x"ffffff",
   21841 => x"fffeb0",
   21842 => x"c30c30",
   21843 => x"c30c30",
   21844 => x"c30c30",
   21845 => x"c30c30",
   21846 => x"c30c30",
   21847 => x"c30c30",
   21848 => x"c30c30",
   21849 => x"c30c30",
   21850 => x"c30c30",
   21851 => x"c30c30",
   21852 => x"c30c30",
   21853 => x"820820",
   21854 => x"820820",
   21855 => x"820820",
   21856 => x"820820",
   21857 => x"820820",
   21858 => x"820820",
   21859 => x"820820",
   21860 => x"820820",
   21861 => x"820820",
   21862 => x"820820",
   21863 => x"820820",
   21864 => x"820820",
   21865 => x"820820",
   21866 => x"820820",
   21867 => x"820820",
   21868 => x"820820",
   21869 => x"820820",
   21870 => x"820820",
   21871 => x"820820",
   21872 => x"820820",
   21873 => x"820820",
   21874 => x"820820",
   21875 => x"820410",
   21876 => x"410410",
   21877 => x"410410",
   21878 => x"410410",
   21879 => x"410410",
   21880 => x"410410",
   21881 => x"410410",
   21882 => x"410410",
   21883 => x"410410",
   21884 => x"410410",
   21885 => x"410410",
   21886 => x"410410",
   21887 => x"410410",
   21888 => x"410410",
   21889 => x"410410",
   21890 => x"410410",
   21891 => x"410410",
   21892 => x"410410",
   21893 => x"410410",
   21894 => x"410410",
   21895 => x"410410",
   21896 => x"410410",
   21897 => x"410410",
   21898 => x"410000",
   21899 => x"000000",
   21900 => x"000000",
   21901 => x"000000",
   21902 => x"000000",
   21903 => x"000000",
   21904 => x"000000",
   21905 => x"000000",
   21906 => x"000000",
   21907 => x"000000",
   21908 => x"000000",
   21909 => x"00057f",
   21910 => x"ffffff",
   21911 => x"ffffff",
   21912 => x"ffffff",
   21913 => x"ffffff",
   21914 => x"ffffff",
   21915 => x"ffffff",
   21916 => x"ffffff",
   21917 => x"ffffff",
   21918 => x"ffffff",
   21919 => x"ffffff",
   21920 => x"ffffff",
   21921 => x"fffff5",
   21922 => x"c30c30",
   21923 => x"c30c30",
   21924 => x"c30c30",
   21925 => x"c30c30",
   21926 => x"c30c30",
   21927 => x"c30c30",
   21928 => x"c30c30",
   21929 => x"c30c30",
   21930 => x"c30c30",
   21931 => x"c30c30",
   21932 => x"c30c30",
   21933 => x"c30c30",
   21934 => x"c30c30",
   21935 => x"c30867",
   21936 => x"df3cf3",
   21937 => x"cf3cf3",
   21938 => x"cf3cf3",
   21939 => x"cf3cf3",
   21940 => x"cf3cf3",
   21941 => x"cf3cf3",
   21942 => x"cf3cf3",
   21943 => x"cf3aae",
   21944 => x"ffffff",
   21945 => x"ffffff",
   21946 => x"ffffff",
   21947 => x"ffffff",
   21948 => x"ffffff",
   21949 => x"ffffff",
   21950 => x"ffffff",
   21951 => x"ffffff",
   21952 => x"ffffff",
   21953 => x"ffffff",
   21954 => x"ffffff",
   21955 => x"ffffff",
   21956 => x"ffffff",
   21957 => x"ffffff",
   21958 => x"ffffff",
   21959 => x"ffffff",
   21960 => x"ffffff",
   21961 => x"ffffff",
   21962 => x"ffffff",
   21963 => x"ffffff",
   21964 => x"ffffde",
   21965 => x"38f3cf",
   21966 => x"3cf3cf",
   21967 => x"3cf3cf",
   21968 => x"3cf3cf",
   21969 => x"3cf3cf",
   21970 => x"3cf3cf",
   21971 => x"3cf3cf",
   21972 => x"3cf3cd",
   21973 => x"30c30c",
   21974 => x"30c30c",
   21975 => x"30c30c",
   21976 => x"30c30c",
   21977 => x"30c30c",
   21978 => x"30c30c",
   21979 => x"30c30c",
   21980 => x"30c30c",
   21981 => x"30c30c",
   21982 => x"30c30c",
   21983 => x"30c30c",
   21984 => x"30c30c",
   21985 => x"30c30c",
   21986 => x"30c32e",
   21987 => x"ffffff",
   21988 => x"ffffff",
   21989 => x"ffffff",
   21990 => x"ffffff",
   21991 => x"ffffff",
   21992 => x"ffffff",
   21993 => x"ffffff",
   21994 => x"ffffff",
   21995 => x"ffffff",
   21996 => x"ffffff",
   21997 => x"fea56a",
   21998 => x"ffffff",
   21999 => x"ffffff",
   22000 => x"ffffff",
   22001 => x"fffeb0",
   22002 => x"c30c30",
   22003 => x"c30c30",
   22004 => x"c30c30",
   22005 => x"c30c30",
   22006 => x"c30c30",
   22007 => x"c30c30",
   22008 => x"c30c30",
   22009 => x"c30c30",
   22010 => x"c30c30",
   22011 => x"c30c30",
   22012 => x"c30c30",
   22013 => x"820820",
   22014 => x"820820",
   22015 => x"820820",
   22016 => x"820820",
   22017 => x"820820",
   22018 => x"820820",
   22019 => x"820820",
   22020 => x"820820",
   22021 => x"820820",
   22022 => x"820820",
   22023 => x"820820",
   22024 => x"820820",
   22025 => x"820820",
   22026 => x"820820",
   22027 => x"820820",
   22028 => x"820820",
   22029 => x"820820",
   22030 => x"820820",
   22031 => x"820820",
   22032 => x"820820",
   22033 => x"820820",
   22034 => x"820820",
   22035 => x"820410",
   22036 => x"410410",
   22037 => x"410410",
   22038 => x"410410",
   22039 => x"410410",
   22040 => x"410410",
   22041 => x"410410",
   22042 => x"410410",
   22043 => x"410410",
   22044 => x"410410",
   22045 => x"410410",
   22046 => x"410410",
   22047 => x"410410",
   22048 => x"410410",
   22049 => x"410410",
   22050 => x"410410",
   22051 => x"410410",
   22052 => x"410410",
   22053 => x"410410",
   22054 => x"410410",
   22055 => x"410410",
   22056 => x"410410",
   22057 => x"410410",
   22058 => x"410000",
   22059 => x"000000",
   22060 => x"000000",
   22061 => x"000000",
   22062 => x"000000",
   22063 => x"000000",
   22064 => x"000000",
   22065 => x"000000",
   22066 => x"000000",
   22067 => x"000000",
   22068 => x"000000",
   22069 => x"00057f",
   22070 => x"ffffff",
   22071 => x"ffffff",
   22072 => x"ffffff",
   22073 => x"ffffff",
   22074 => x"ffffff",
   22075 => x"ffffff",
   22076 => x"ffffff",
   22077 => x"ffffff",
   22078 => x"ffffff",
   22079 => x"ffffff",
   22080 => x"ffffff",
   22081 => x"fffffa",
   22082 => x"c30c30",
   22083 => x"c30c30",
   22084 => x"c30c30",
   22085 => x"c30c30",
   22086 => x"c30c30",
   22087 => x"c30c30",
   22088 => x"c30c30",
   22089 => x"c30c30",
   22090 => x"c30c30",
   22091 => x"c30c30",
   22092 => x"c30c30",
   22093 => x"c30c30",
   22094 => x"c30c30",
   22095 => x"c219b7",
   22096 => x"cf3cf3",
   22097 => x"cf3cf3",
   22098 => x"cf3cf3",
   22099 => x"cf3cf3",
   22100 => x"cf3cf3",
   22101 => x"cf3cf3",
   22102 => x"cf3cf3",
   22103 => x"cf39aa",
   22104 => x"ffffff",
   22105 => x"ffffff",
   22106 => x"ffffff",
   22107 => x"ffffff",
   22108 => x"ffffff",
   22109 => x"ffffff",
   22110 => x"ffffff",
   22111 => x"ffffff",
   22112 => x"ffffff",
   22113 => x"ffffff",
   22114 => x"ffffff",
   22115 => x"ffffff",
   22116 => x"ffffff",
   22117 => x"ffffff",
   22118 => x"ffffff",
   22119 => x"ffffff",
   22120 => x"ffffff",
   22121 => x"ffffff",
   22122 => x"ffffff",
   22123 => x"ffffff",
   22124 => x"fffb9d",
   22125 => x"3cf3cf",
   22126 => x"3cf3cf",
   22127 => x"3cf3cf",
   22128 => x"3cf3cf",
   22129 => x"3cf3cf",
   22130 => x"3cf3cf",
   22131 => x"3cf3cf",
   22132 => x"3cf3ce",
   22133 => x"30c30c",
   22134 => x"30c30c",
   22135 => x"30c30c",
   22136 => x"30c30c",
   22137 => x"30c30c",
   22138 => x"30c30c",
   22139 => x"30c30c",
   22140 => x"30c30c",
   22141 => x"30c30c",
   22142 => x"30c30c",
   22143 => x"30c30c",
   22144 => x"30c30c",
   22145 => x"30c30c",
   22146 => x"30c77f",
   22147 => x"ffffff",
   22148 => x"ffffff",
   22149 => x"ffffff",
   22150 => x"ffffff",
   22151 => x"ffffff",
   22152 => x"ffffff",
   22153 => x"ffffff",
   22154 => x"ffffff",
   22155 => x"ffffff",
   22156 => x"ffffff",
   22157 => x"a95abf",
   22158 => x"ffffff",
   22159 => x"ffffff",
   22160 => x"ffffff",
   22161 => x"fffeb0",
   22162 => x"c30c30",
   22163 => x"c30c30",
   22164 => x"c30c30",
   22165 => x"c30c30",
   22166 => x"c30c30",
   22167 => x"c30c30",
   22168 => x"c30c30",
   22169 => x"c30c30",
   22170 => x"c30c30",
   22171 => x"c30c30",
   22172 => x"c30c30",
   22173 => x"820820",
   22174 => x"820820",
   22175 => x"820820",
   22176 => x"820820",
   22177 => x"820820",
   22178 => x"820820",
   22179 => x"820820",
   22180 => x"820820",
   22181 => x"820820",
   22182 => x"820820",
   22183 => x"820820",
   22184 => x"820820",
   22185 => x"820820",
   22186 => x"820820",
   22187 => x"820820",
   22188 => x"820820",
   22189 => x"820820",
   22190 => x"820820",
   22191 => x"820820",
   22192 => x"820820",
   22193 => x"820820",
   22194 => x"820820",
   22195 => x"820410",
   22196 => x"410410",
   22197 => x"410410",
   22198 => x"410410",
   22199 => x"410410",
   22200 => x"410410",
   22201 => x"410410",
   22202 => x"410410",
   22203 => x"410410",
   22204 => x"410410",
   22205 => x"410410",
   22206 => x"410410",
   22207 => x"410410",
   22208 => x"410410",
   22209 => x"410410",
   22210 => x"410410",
   22211 => x"410410",
   22212 => x"410410",
   22213 => x"410410",
   22214 => x"410410",
   22215 => x"410410",
   22216 => x"410410",
   22217 => x"410410",
   22218 => x"410000",
   22219 => x"000000",
   22220 => x"000000",
   22221 => x"000000",
   22222 => x"000000",
   22223 => x"000000",
   22224 => x"000000",
   22225 => x"000000",
   22226 => x"000000",
   22227 => x"000000",
   22228 => x"000000",
   22229 => x"00057f",
   22230 => x"ffffff",
   22231 => x"ffffff",
   22232 => x"ffffff",
   22233 => x"ffffff",
   22234 => x"ffffff",
   22235 => x"ffffff",
   22236 => x"ffffff",
   22237 => x"ffffff",
   22238 => x"ffffff",
   22239 => x"ffffff",
   22240 => x"ffffff",
   22241 => x"ffffff",
   22242 => x"d70c30",
   22243 => x"c30c30",
   22244 => x"c30c30",
   22245 => x"c30c30",
   22246 => x"c30c30",
   22247 => x"c30c30",
   22248 => x"c30c30",
   22249 => x"c30c30",
   22250 => x"c30c30",
   22251 => x"c30c30",
   22252 => x"c30c30",
   22253 => x"c30c30",
   22254 => x"c30c30",
   22255 => x"8269f3",
   22256 => x"cf3cf3",
   22257 => x"cf3cf3",
   22258 => x"cf3cf3",
   22259 => x"cf3cf3",
   22260 => x"cf3cf3",
   22261 => x"cf3cf3",
   22262 => x"cf3cf3",
   22263 => x"cf3cea",
   22264 => x"bbffff",
   22265 => x"ffffff",
   22266 => x"ffffff",
   22267 => x"ffffff",
   22268 => x"ffffff",
   22269 => x"ffffff",
   22270 => x"ffffff",
   22271 => x"ffffff",
   22272 => x"ffffff",
   22273 => x"ffffff",
   22274 => x"ffffff",
   22275 => x"ffffff",
   22276 => x"ffffff",
   22277 => x"ffffff",
   22278 => x"ffffff",
   22279 => x"ffffff",
   22280 => x"ffffff",
   22281 => x"ffffff",
   22282 => x"ffffff",
   22283 => x"ffffff",
   22284 => x"fffb8e",
   22285 => x"3cf3cf",
   22286 => x"3cf3cf",
   22287 => x"3cf3cf",
   22288 => x"3cf3cf",
   22289 => x"3cf3cf",
   22290 => x"3cf3cf",
   22291 => x"3cf3cf",
   22292 => x"3cf3cf",
   22293 => x"38c30c",
   22294 => x"30c30c",
   22295 => x"30c30c",
   22296 => x"30c30c",
   22297 => x"30c30c",
   22298 => x"30c30c",
   22299 => x"30c30c",
   22300 => x"30c30c",
   22301 => x"30c30c",
   22302 => x"30c30c",
   22303 => x"30c30c",
   22304 => x"30c30c",
   22305 => x"30c30c",
   22306 => x"30cbbf",
   22307 => x"ffffff",
   22308 => x"ffffff",
   22309 => x"ffffff",
   22310 => x"ffffff",
   22311 => x"ffffff",
   22312 => x"ffffff",
   22313 => x"ffffff",
   22314 => x"ffffff",
   22315 => x"ffffff",
   22316 => x"ffffea",
   22317 => x"56afff",
   22318 => x"ffffff",
   22319 => x"ffffff",
   22320 => x"ffffff",
   22321 => x"fffeb0",
   22322 => x"c30c30",
   22323 => x"c30c30",
   22324 => x"c30c30",
   22325 => x"c30c30",
   22326 => x"c30c30",
   22327 => x"c30c30",
   22328 => x"c30c30",
   22329 => x"c30c30",
   22330 => x"c30c30",
   22331 => x"c30c30",
   22332 => x"c30c30",
   22333 => x"820820",
   22334 => x"820820",
   22335 => x"820820",
   22336 => x"820820",
   22337 => x"820820",
   22338 => x"820820",
   22339 => x"820820",
   22340 => x"820820",
   22341 => x"820820",
   22342 => x"820820",
   22343 => x"820820",
   22344 => x"820820",
   22345 => x"820820",
   22346 => x"820820",
   22347 => x"820820",
   22348 => x"820820",
   22349 => x"820820",
   22350 => x"820820",
   22351 => x"820820",
   22352 => x"820820",
   22353 => x"820820",
   22354 => x"820820",
   22355 => x"820410",
   22356 => x"410410",
   22357 => x"410410",
   22358 => x"410410",
   22359 => x"410410",
   22360 => x"410410",
   22361 => x"410410",
   22362 => x"410410",
   22363 => x"410410",
   22364 => x"410410",
   22365 => x"410410",
   22366 => x"410410",
   22367 => x"410410",
   22368 => x"410410",
   22369 => x"410410",
   22370 => x"410410",
   22371 => x"410410",
   22372 => x"410410",
   22373 => x"410410",
   22374 => x"410410",
   22375 => x"410410",
   22376 => x"410410",
   22377 => x"410410",
   22378 => x"410000",
   22379 => x"000000",
   22380 => x"000000",
   22381 => x"000000",
   22382 => x"000000",
   22383 => x"000000",
   22384 => x"000000",
   22385 => x"000000",
   22386 => x"000000",
   22387 => x"000000",
   22388 => x"000000",
   22389 => x"00057f",
   22390 => x"ffffff",
   22391 => x"ffffff",
   22392 => x"ffffff",
   22393 => x"ffffff",
   22394 => x"ffffff",
   22395 => x"ffffff",
   22396 => x"ffffff",
   22397 => x"ffffff",
   22398 => x"ffffff",
   22399 => x"ffffff",
   22400 => x"ffffff",
   22401 => x"ffffff",
   22402 => x"d70c30",
   22403 => x"c30c30",
   22404 => x"c30c30",
   22405 => x"c30c30",
   22406 => x"c30c30",
   22407 => x"c30c30",
   22408 => x"c30c30",
   22409 => x"c30c30",
   22410 => x"c30c30",
   22411 => x"c30c30",
   22412 => x"c30c30",
   22413 => x"c30c30",
   22414 => x"c30c30",
   22415 => x"8a7df3",
   22416 => x"cf3cf3",
   22417 => x"cf3cf3",
   22418 => x"cf3cf3",
   22419 => x"cf3cf3",
   22420 => x"cf3cf3",
   22421 => x"cf3cf3",
   22422 => x"cf3cf3",
   22423 => x"cf3ce6",
   22424 => x"bbffff",
   22425 => x"ffffff",
   22426 => x"ffffff",
   22427 => x"ffffff",
   22428 => x"ffffff",
   22429 => x"ffffff",
   22430 => x"ffffff",
   22431 => x"ffffff",
   22432 => x"ffffff",
   22433 => x"ffffff",
   22434 => x"ffffff",
   22435 => x"ffffff",
   22436 => x"ffffff",
   22437 => x"ffffff",
   22438 => x"ffffff",
   22439 => x"ffffff",
   22440 => x"ffffff",
   22441 => x"ffffff",
   22442 => x"ffffff",
   22443 => x"ffffff",
   22444 => x"fff78e",
   22445 => x"3cf3cf",
   22446 => x"3cf3cf",
   22447 => x"3cf3cf",
   22448 => x"3cf3cf",
   22449 => x"3cf3cf",
   22450 => x"3cf3cf",
   22451 => x"3cf3cf",
   22452 => x"3cf3cf",
   22453 => x"3cd30c",
   22454 => x"30c30c",
   22455 => x"30c30c",
   22456 => x"30c30c",
   22457 => x"30c30c",
   22458 => x"30c30c",
   22459 => x"30c30c",
   22460 => x"30c30c",
   22461 => x"30c30c",
   22462 => x"30c30c",
   22463 => x"30c30c",
   22464 => x"30c30c",
   22465 => x"30c30c",
   22466 => x"30cbbf",
   22467 => x"ffffff",
   22468 => x"ffffff",
   22469 => x"ffffff",
   22470 => x"ffffff",
   22471 => x"ffffff",
   22472 => x"ffffff",
   22473 => x"ffffff",
   22474 => x"ffffff",
   22475 => x"ffffff",
   22476 => x"fffa95",
   22477 => x"abffff",
   22478 => x"ffffff",
   22479 => x"ffffff",
   22480 => x"ffffff",
   22481 => x"fffeb0",
   22482 => x"c30c30",
   22483 => x"c30c30",
   22484 => x"c30c30",
   22485 => x"c30c30",
   22486 => x"c30c30",
   22487 => x"c30c30",
   22488 => x"c30c30",
   22489 => x"c30c30",
   22490 => x"c30c30",
   22491 => x"c30c30",
   22492 => x"c30c30",
   22493 => x"820820",
   22494 => x"820820",
   22495 => x"820820",
   22496 => x"820820",
   22497 => x"820820",
   22498 => x"820820",
   22499 => x"820820",
   22500 => x"820820",
   22501 => x"820820",
   22502 => x"820820",
   22503 => x"820820",
   22504 => x"820820",
   22505 => x"820820",
   22506 => x"820820",
   22507 => x"820820",
   22508 => x"820820",
   22509 => x"820820",
   22510 => x"820820",
   22511 => x"820820",
   22512 => x"820820",
   22513 => x"820820",
   22514 => x"820820",
   22515 => x"820410",
   22516 => x"410410",
   22517 => x"410410",
   22518 => x"410410",
   22519 => x"410410",
   22520 => x"410410",
   22521 => x"410410",
   22522 => x"410410",
   22523 => x"410410",
   22524 => x"410410",
   22525 => x"410410",
   22526 => x"410410",
   22527 => x"410410",
   22528 => x"410410",
   22529 => x"410410",
   22530 => x"410410",
   22531 => x"410410",
   22532 => x"410410",
   22533 => x"410410",
   22534 => x"410410",
   22535 => x"410410",
   22536 => x"410410",
   22537 => x"410410",
   22538 => x"410000",
   22539 => x"000000",
   22540 => x"000000",
   22541 => x"000000",
   22542 => x"000000",
   22543 => x"000000",
   22544 => x"000000",
   22545 => x"000000",
   22546 => x"000000",
   22547 => x"000000",
   22548 => x"000000",
   22549 => x"00057f",
   22550 => x"ffffff",
   22551 => x"ffffff",
   22552 => x"ffffff",
   22553 => x"ffffff",
   22554 => x"ffffff",
   22555 => x"ffffff",
   22556 => x"ffffff",
   22557 => x"ffffff",
   22558 => x"ffffff",
   22559 => x"ffffff",
   22560 => x"ffffff",
   22561 => x"ffffff",
   22562 => x"eb5c30",
   22563 => x"c30c30",
   22564 => x"c30c30",
   22565 => x"c30c30",
   22566 => x"c30c30",
   22567 => x"c30c30",
   22568 => x"c30c30",
   22569 => x"c30c30",
   22570 => x"c30c30",
   22571 => x"c30c30",
   22572 => x"c30c30",
   22573 => x"c30c30",
   22574 => x"c30c21",
   22575 => x"9f7cf3",
   22576 => x"cf3cf3",
   22577 => x"cf3cf3",
   22578 => x"cf3cf3",
   22579 => x"cf3cf3",
   22580 => x"cf3cf3",
   22581 => x"cf3cf3",
   22582 => x"cf3cf3",
   22583 => x"cf3cf7",
   22584 => x"abffff",
   22585 => x"ffffff",
   22586 => x"ffffff",
   22587 => x"ffffff",
   22588 => x"ffffff",
   22589 => x"ffffff",
   22590 => x"ffffff",
   22591 => x"ffffff",
   22592 => x"ffffff",
   22593 => x"ffffff",
   22594 => x"ffffff",
   22595 => x"ffffff",
   22596 => x"ffffff",
   22597 => x"ffffff",
   22598 => x"ffffff",
   22599 => x"ffffff",
   22600 => x"ffffff",
   22601 => x"ffffff",
   22602 => x"ffffff",
   22603 => x"ffffff",
   22604 => x"fee38f",
   22605 => x"3cf3cf",
   22606 => x"3cf3cf",
   22607 => x"3cf3cf",
   22608 => x"3cf3cf",
   22609 => x"3cf3cf",
   22610 => x"3cf3cf",
   22611 => x"3cf3cf",
   22612 => x"3cf3cf",
   22613 => x"3ce34c",
   22614 => x"30c30c",
   22615 => x"30c30c",
   22616 => x"30c30c",
   22617 => x"30c30c",
   22618 => x"30c30c",
   22619 => x"30c30c",
   22620 => x"30c30c",
   22621 => x"30c30c",
   22622 => x"30c30c",
   22623 => x"30c30c",
   22624 => x"30c30c",
   22625 => x"30c30c",
   22626 => x"31dfff",
   22627 => x"ffffff",
   22628 => x"ffffff",
   22629 => x"ffffff",
   22630 => x"ffffff",
   22631 => x"ffffff",
   22632 => x"ffffff",
   22633 => x"ffffff",
   22634 => x"ffffff",
   22635 => x"ffffff",
   22636 => x"fea56a",
   22637 => x"ffffff",
   22638 => x"ffffff",
   22639 => x"ffffff",
   22640 => x"ffffff",
   22641 => x"fffeb0",
   22642 => x"c30c30",
   22643 => x"c30c30",
   22644 => x"c30c30",
   22645 => x"c30c30",
   22646 => x"c30c30",
   22647 => x"c30c30",
   22648 => x"c30c30",
   22649 => x"c30c30",
   22650 => x"c30c30",
   22651 => x"c30c30",
   22652 => x"c30c30",
   22653 => x"820820",
   22654 => x"820820",
   22655 => x"820820",
   22656 => x"820820",
   22657 => x"820820",
   22658 => x"820820",
   22659 => x"820820",
   22660 => x"820820",
   22661 => x"820820",
   22662 => x"820820",
   22663 => x"820820",
   22664 => x"820820",
   22665 => x"820820",
   22666 => x"820820",
   22667 => x"820820",
   22668 => x"820820",
   22669 => x"820820",
   22670 => x"820820",
   22671 => x"820820",
   22672 => x"820820",
   22673 => x"820820",
   22674 => x"820820",
   22675 => x"820410",
   22676 => x"410410",
   22677 => x"410410",
   22678 => x"410410",
   22679 => x"410410",
   22680 => x"410410",
   22681 => x"410410",
   22682 => x"410410",
   22683 => x"410410",
   22684 => x"410410",
   22685 => x"410410",
   22686 => x"410410",
   22687 => x"410410",
   22688 => x"410410",
   22689 => x"410410",
   22690 => x"410410",
   22691 => x"410410",
   22692 => x"410410",
   22693 => x"410410",
   22694 => x"410410",
   22695 => x"410410",
   22696 => x"410410",
   22697 => x"410410",
   22698 => x"410000",
   22699 => x"000000",
   22700 => x"000000",
   22701 => x"000000",
   22702 => x"000000",
   22703 => x"000000",
   22704 => x"000000",
   22705 => x"000000",
   22706 => x"000000",
   22707 => x"000000",
   22708 => x"000000",
   22709 => x"00057f",
   22710 => x"ffffff",
   22711 => x"ffffff",
   22712 => x"ffffff",
   22713 => x"ffffea",
   22714 => x"aaaaaa",
   22715 => x"aaaaaa",
   22716 => x"aaaaaa",
   22717 => x"ffffff",
   22718 => x"ffffff",
   22719 => x"ffffff",
   22720 => x"ffffff",
   22721 => x"ffffff",
   22722 => x"ff5c30",
   22723 => x"c30c30",
   22724 => x"c30c30",
   22725 => x"c30c30",
   22726 => x"c30c30",
   22727 => x"c30c30",
   22728 => x"c30c30",
   22729 => x"c30c30",
   22730 => x"c30c30",
   22731 => x"c30c30",
   22732 => x"c30c30",
   22733 => x"c30c30",
   22734 => x"c30c16",
   22735 => x"9f3cf3",
   22736 => x"cf3cf3",
   22737 => x"cf3cf3",
   22738 => x"cf3cf3",
   22739 => x"cf3cf3",
   22740 => x"cf3cf3",
   22741 => x"cf3cf3",
   22742 => x"cf3cf3",
   22743 => x"cf3cf3",
   22744 => x"9aefff",
   22745 => x"ffffff",
   22746 => x"ffffff",
   22747 => x"ffffff",
   22748 => x"ffffff",
   22749 => x"ffffff",
   22750 => x"ffffff",
   22751 => x"ffffff",
   22752 => x"ffffff",
   22753 => x"ffffff",
   22754 => x"ffffff",
   22755 => x"ffffff",
   22756 => x"ffffff",
   22757 => x"ffffff",
   22758 => x"ffffff",
   22759 => x"ffffff",
   22760 => x"ffffff",
   22761 => x"ffffff",
   22762 => x"ffffff",
   22763 => x"ffffff",
   22764 => x"fee38f",
   22765 => x"3cf3cf",
   22766 => x"3cf3cf",
   22767 => x"3cf3cf",
   22768 => x"3cf3cf",
   22769 => x"3cf3cf",
   22770 => x"3cf3cf",
   22771 => x"3cf3cf",
   22772 => x"3cf3cf",
   22773 => x"3cf38c",
   22774 => x"30c30c",
   22775 => x"30c30c",
   22776 => x"30c30c",
   22777 => x"30c30c",
   22778 => x"30c30c",
   22779 => x"30c30c",
   22780 => x"30c30c",
   22781 => x"30c30c",
   22782 => x"30c30c",
   22783 => x"30c30c",
   22784 => x"30c30c",
   22785 => x"30c30c",
   22786 => x"32efff",
   22787 => x"ffffff",
   22788 => x"ffffff",
   22789 => x"ffffff",
   22790 => x"ffffff",
   22791 => x"ffffff",
   22792 => x"ffffff",
   22793 => x"ffffff",
   22794 => x"ffffff",
   22795 => x"ffffff",
   22796 => x"a95abf",
   22797 => x"ffffff",
   22798 => x"ffffff",
   22799 => x"ffffff",
   22800 => x"ffffff",
   22801 => x"fffeb0",
   22802 => x"c30c30",
   22803 => x"c30c30",
   22804 => x"c30c30",
   22805 => x"c30c30",
   22806 => x"c30c30",
   22807 => x"c30c30",
   22808 => x"c30c30",
   22809 => x"c30c30",
   22810 => x"c30c30",
   22811 => x"c30c30",
   22812 => x"c30c30",
   22813 => x"820820",
   22814 => x"820820",
   22815 => x"820820",
   22816 => x"820820",
   22817 => x"820820",
   22818 => x"820820",
   22819 => x"820820",
   22820 => x"820820",
   22821 => x"820820",
   22822 => x"820820",
   22823 => x"820820",
   22824 => x"820820",
   22825 => x"820820",
   22826 => x"820820",
   22827 => x"820820",
   22828 => x"820820",
   22829 => x"820820",
   22830 => x"820820",
   22831 => x"820820",
   22832 => x"820820",
   22833 => x"820820",
   22834 => x"820820",
   22835 => x"820410",
   22836 => x"410410",
   22837 => x"410410",
   22838 => x"410410",
   22839 => x"410410",
   22840 => x"410410",
   22841 => x"410410",
   22842 => x"410410",
   22843 => x"410410",
   22844 => x"410410",
   22845 => x"410410",
   22846 => x"410410",
   22847 => x"410410",
   22848 => x"410410",
   22849 => x"410410",
   22850 => x"410410",
   22851 => x"410410",
   22852 => x"410410",
   22853 => x"410410",
   22854 => x"410410",
   22855 => x"410410",
   22856 => x"410410",
   22857 => x"410410",
   22858 => x"410000",
   22859 => x"000000",
   22860 => x"000000",
   22861 => x"000000",
   22862 => x"000000",
   22863 => x"000000",
   22864 => x"000000",
   22865 => x"000000",
   22866 => x"000000",
   22867 => x"000000",
   22868 => x"000000",
   22869 => x"00057f",
   22870 => x"ffffff",
   22871 => x"ffffff",
   22872 => x"ffffff",
   22873 => x"ffffd5",
   22874 => x"000000",
   22875 => x"000000",
   22876 => x"000015",
   22877 => x"555abf",
   22878 => x"ffffff",
   22879 => x"ffffff",
   22880 => x"ffffff",
   22881 => x"ffffff",
   22882 => x"ffad70",
   22883 => x"c30c30",
   22884 => x"c30c30",
   22885 => x"c30c30",
   22886 => x"c30c30",
   22887 => x"c30c30",
   22888 => x"c30c30",
   22889 => x"c30c30",
   22890 => x"c30c30",
   22891 => x"c30c30",
   22892 => x"c30c30",
   22893 => x"c30c30",
   22894 => x"c30867",
   22895 => x"cf3cf3",
   22896 => x"cf3cf3",
   22897 => x"cf3cf3",
   22898 => x"cf3cf3",
   22899 => x"cf3cf3",
   22900 => x"cf3cf3",
   22901 => x"cf3cf3",
   22902 => x"cf3cf3",
   22903 => x"cf3cf3",
   22904 => x"9eafff",
   22905 => x"ffffff",
   22906 => x"ffffff",
   22907 => x"ffffff",
   22908 => x"ffffff",
   22909 => x"ffffff",
   22910 => x"ffffff",
   22911 => x"ffffff",
   22912 => x"ffffff",
   22913 => x"ffffff",
   22914 => x"ffffff",
   22915 => x"ffffff",
   22916 => x"ffffff",
   22917 => x"ffffff",
   22918 => x"ffffff",
   22919 => x"ffffff",
   22920 => x"ffffff",
   22921 => x"ffffff",
   22922 => x"ffffff",
   22923 => x"ffffff",
   22924 => x"b9e3cf",
   22925 => x"3cf3cf",
   22926 => x"3cf3cf",
   22927 => x"3cf3cf",
   22928 => x"3cf3cf",
   22929 => x"3cf3cf",
   22930 => x"3cf3cf",
   22931 => x"3cf3cf",
   22932 => x"3cf3cf",
   22933 => x"3cf3cd",
   22934 => x"30c30c",
   22935 => x"30c30c",
   22936 => x"30c30c",
   22937 => x"30c30c",
   22938 => x"30c30c",
   22939 => x"30c30c",
   22940 => x"30c30c",
   22941 => x"30c30c",
   22942 => x"30c30c",
   22943 => x"30c30c",
   22944 => x"30c30c",
   22945 => x"30c30c",
   22946 => x"77ffff",
   22947 => x"ffffff",
   22948 => x"ffffff",
   22949 => x"ffffff",
   22950 => x"ffffff",
   22951 => x"ffffff",
   22952 => x"ffffff",
   22953 => x"ffffff",
   22954 => x"ffffff",
   22955 => x"ffffea",
   22956 => x"56afff",
   22957 => x"ffffff",
   22958 => x"ffffff",
   22959 => x"ffffff",
   22960 => x"ffffff",
   22961 => x"fffeb0",
   22962 => x"c30c30",
   22963 => x"c30c30",
   22964 => x"c30c30",
   22965 => x"c30c30",
   22966 => x"c30c30",
   22967 => x"c30c30",
   22968 => x"c30c30",
   22969 => x"c30c30",
   22970 => x"c30c30",
   22971 => x"c30c30",
   22972 => x"c30c30",
   22973 => x"820820",
   22974 => x"820820",
   22975 => x"820820",
   22976 => x"820820",
   22977 => x"820820",
   22978 => x"820820",
   22979 => x"820820",
   22980 => x"820820",
   22981 => x"820820",
   22982 => x"820820",
   22983 => x"820820",
   22984 => x"820820",
   22985 => x"820820",
   22986 => x"820820",
   22987 => x"820820",
   22988 => x"820820",
   22989 => x"820820",
   22990 => x"820820",
   22991 => x"820820",
   22992 => x"820820",
   22993 => x"820820",
   22994 => x"820820",
   22995 => x"820410",
   22996 => x"410410",
   22997 => x"410410",
   22998 => x"410410",
   22999 => x"410410",
   23000 => x"410410",
   23001 => x"410410",
   23002 => x"410410",
   23003 => x"410410",
   23004 => x"410410",
   23005 => x"410410",
   23006 => x"410410",
   23007 => x"410410",
   23008 => x"410410",
   23009 => x"410410",
   23010 => x"410410",
   23011 => x"410410",
   23012 => x"410410",
   23013 => x"410410",
   23014 => x"410410",
   23015 => x"410410",
   23016 => x"410410",
   23017 => x"410410",
   23018 => x"410000",
   23019 => x"000000",
   23020 => x"000000",
   23021 => x"000000",
   23022 => x"000000",
   23023 => x"000000",
   23024 => x"000000",
   23025 => x"000000",
   23026 => x"000000",
   23027 => x"000000",
   23028 => x"000000",
   23029 => x"00057f",
   23030 => x"ffffff",
   23031 => x"ffffff",
   23032 => x"ffffff",
   23033 => x"ffffd5",
   23034 => x"000000",
   23035 => x"000000",
   23036 => x"000000",
   23037 => x"000015",
   23038 => x"abffff",
   23039 => x"ffffff",
   23040 => x"ffffff",
   23041 => x"ffffff",
   23042 => x"fffd70",
   23043 => x"c30c30",
   23044 => x"c30c30",
   23045 => x"c30c30",
   23046 => x"c30c30",
   23047 => x"c30c30",
   23048 => x"c30c30",
   23049 => x"c30c30",
   23050 => x"c30c30",
   23051 => x"c30c30",
   23052 => x"c30c30",
   23053 => x"c30c30",
   23054 => x"c215b7",
   23055 => x"cf3cf3",
   23056 => x"cf3cf3",
   23057 => x"cf3cf3",
   23058 => x"cf3cf3",
   23059 => x"cf3cf3",
   23060 => x"cf3cf3",
   23061 => x"cf3cf3",
   23062 => x"cf3cf3",
   23063 => x"cf3cf3",
   23064 => x"ceabbf",
   23065 => x"ffffff",
   23066 => x"ffffff",
   23067 => x"ffffff",
   23068 => x"ffffff",
   23069 => x"ffffff",
   23070 => x"ffffff",
   23071 => x"ffffff",
   23072 => x"ffffff",
   23073 => x"ffffff",
   23074 => x"ffffff",
   23075 => x"ffffff",
   23076 => x"ffffff",
   23077 => x"ffffff",
   23078 => x"ffffff",
   23079 => x"ffffff",
   23080 => x"ffffff",
   23081 => x"ffffff",
   23082 => x"ffffff",
   23083 => x"ffffff",
   23084 => x"b8e3cf",
   23085 => x"3cf3cf",
   23086 => x"3cf3cf",
   23087 => x"3cf3cf",
   23088 => x"3cf3cf",
   23089 => x"3cf3cf",
   23090 => x"3cf3cf",
   23091 => x"3cf3cf",
   23092 => x"3cf3cf",
   23093 => x"3cf3ce",
   23094 => x"30c30c",
   23095 => x"30c30c",
   23096 => x"30c30c",
   23097 => x"30c30c",
   23098 => x"30c30c",
   23099 => x"30c30c",
   23100 => x"30c30c",
   23101 => x"30c30c",
   23102 => x"30c30c",
   23103 => x"30c30c",
   23104 => x"30c30c",
   23105 => x"30c30c",
   23106 => x"bbffff",
   23107 => x"ffffff",
   23108 => x"ffffff",
   23109 => x"ffffff",
   23110 => x"ffffff",
   23111 => x"ffffff",
   23112 => x"ffffff",
   23113 => x"ffffff",
   23114 => x"ffffff",
   23115 => x"fffa95",
   23116 => x"abffff",
   23117 => x"ffffff",
   23118 => x"ffffff",
   23119 => x"ffffff",
   23120 => x"ffffff",
   23121 => x"fffeb0",
   23122 => x"c30c30",
   23123 => x"c30c30",
   23124 => x"c30c30",
   23125 => x"c30c30",
   23126 => x"c30c30",
   23127 => x"c30c30",
   23128 => x"c30c30",
   23129 => x"c30c30",
   23130 => x"c30c30",
   23131 => x"c30c30",
   23132 => x"c30c30",
   23133 => x"820820",
   23134 => x"820820",
   23135 => x"820820",
   23136 => x"820820",
   23137 => x"820820",
   23138 => x"820820",
   23139 => x"820820",
   23140 => x"820820",
   23141 => x"820820",
   23142 => x"820820",
   23143 => x"820820",
   23144 => x"820820",
   23145 => x"820820",
   23146 => x"820820",
   23147 => x"820820",
   23148 => x"820820",
   23149 => x"820820",
   23150 => x"820820",
   23151 => x"820820",
   23152 => x"820820",
   23153 => x"820820",
   23154 => x"820820",
   23155 => x"820410",
   23156 => x"410410",
   23157 => x"410410",
   23158 => x"410410",
   23159 => x"410410",
   23160 => x"410410",
   23161 => x"410410",
   23162 => x"410410",
   23163 => x"410410",
   23164 => x"410410",
   23165 => x"410410",
   23166 => x"410410",
   23167 => x"410410",
   23168 => x"410410",
   23169 => x"410410",
   23170 => x"410410",
   23171 => x"410410",
   23172 => x"410410",
   23173 => x"410410",
   23174 => x"410410",
   23175 => x"410410",
   23176 => x"410410",
   23177 => x"410410",
   23178 => x"410000",
   23179 => x"000000",
   23180 => x"000000",
   23181 => x"000000",
   23182 => x"000000",
   23183 => x"000000",
   23184 => x"000000",
   23185 => x"000000",
   23186 => x"000000",
   23187 => x"000000",
   23188 => x"000000",
   23189 => x"00057f",
   23190 => x"ffffff",
   23191 => x"ffffff",
   23192 => x"ffffff",
   23193 => x"ffffd5",
   23194 => x"000000",
   23195 => x"555555",
   23196 => x"540000",
   23197 => x"000000",
   23198 => x"56afff",
   23199 => x"ffffff",
   23200 => x"ffffff",
   23201 => x"ffffff",
   23202 => x"fffeb5",
   23203 => x"c30c30",
   23204 => x"c30c30",
   23205 => x"c30c30",
   23206 => x"c30c30",
   23207 => x"c30c30",
   23208 => x"c30c30",
   23209 => x"c30c30",
   23210 => x"c30c30",
   23211 => x"c30c30",
   23212 => x"c30c30",
   23213 => x"c30c30",
   23214 => x"c129f3",
   23215 => x"cf3cf3",
   23216 => x"cf3cf3",
   23217 => x"cf3cf3",
   23218 => x"cf3cf3",
   23219 => x"cf3cf3",
   23220 => x"cf3cf3",
   23221 => x"cf3cf3",
   23222 => x"cf3cf3",
   23223 => x"cf3cf3",
   23224 => x"ce7abf",
   23225 => x"ffffff",
   23226 => x"ffffff",
   23227 => x"ffffff",
   23228 => x"ffffff",
   23229 => x"ffffff",
   23230 => x"ffffff",
   23231 => x"ffffff",
   23232 => x"ffffff",
   23233 => x"ffffff",
   23234 => x"ffffff",
   23235 => x"ffffff",
   23236 => x"ffffff",
   23237 => x"ffffff",
   23238 => x"ffffff",
   23239 => x"ffffff",
   23240 => x"ffffff",
   23241 => x"ffffff",
   23242 => x"ffffff",
   23243 => x"ffffee",
   23244 => x"78f3cf",
   23245 => x"3cf3cf",
   23246 => x"3cf3cf",
   23247 => x"3cf3cf",
   23248 => x"3cf3cf",
   23249 => x"3cf3cf",
   23250 => x"3cf3cf",
   23251 => x"3cf3cf",
   23252 => x"3cf3cf",
   23253 => x"3cf3cf",
   23254 => x"34c30c",
   23255 => x"30c30c",
   23256 => x"30c30c",
   23257 => x"30c30c",
   23258 => x"30c30c",
   23259 => x"30c30c",
   23260 => x"30c30c",
   23261 => x"30c30c",
   23262 => x"30c30c",
   23263 => x"30c30c",
   23264 => x"30c30c",
   23265 => x"30c31d",
   23266 => x"ffffff",
   23267 => x"ffffff",
   23268 => x"ffffff",
   23269 => x"ffffff",
   23270 => x"ffffff",
   23271 => x"ffffff",
   23272 => x"ffffff",
   23273 => x"ffffff",
   23274 => x"ffffff",
   23275 => x"fea56a",
   23276 => x"ffffff",
   23277 => x"ffffff",
   23278 => x"ffffff",
   23279 => x"ffffff",
   23280 => x"ffffff",
   23281 => x"fffeb0",
   23282 => x"c30c30",
   23283 => x"c30c30",
   23284 => x"c30c30",
   23285 => x"c30c30",
   23286 => x"c30c30",
   23287 => x"c30c30",
   23288 => x"c30c30",
   23289 => x"c30c30",
   23290 => x"c30c30",
   23291 => x"c30c30",
   23292 => x"c30c30",
   23293 => x"820820",
   23294 => x"820820",
   23295 => x"820820",
   23296 => x"820820",
   23297 => x"820820",
   23298 => x"820820",
   23299 => x"820820",
   23300 => x"820820",
   23301 => x"820820",
   23302 => x"820820",
   23303 => x"820820",
   23304 => x"820820",
   23305 => x"820820",
   23306 => x"820820",
   23307 => x"820820",
   23308 => x"820820",
   23309 => x"820820",
   23310 => x"820820",
   23311 => x"820820",
   23312 => x"820820",
   23313 => x"820820",
   23314 => x"820820",
   23315 => x"820410",
   23316 => x"410410",
   23317 => x"410410",
   23318 => x"410410",
   23319 => x"410410",
   23320 => x"410410",
   23321 => x"410410",
   23322 => x"410410",
   23323 => x"410410",
   23324 => x"410410",
   23325 => x"410410",
   23326 => x"410410",
   23327 => x"410410",
   23328 => x"410410",
   23329 => x"410410",
   23330 => x"410410",
   23331 => x"410410",
   23332 => x"410410",
   23333 => x"410410",
   23334 => x"410410",
   23335 => x"410410",
   23336 => x"410410",
   23337 => x"410410",
   23338 => x"410000",
   23339 => x"000000",
   23340 => x"000000",
   23341 => x"000000",
   23342 => x"000000",
   23343 => x"000000",
   23344 => x"000000",
   23345 => x"000000",
   23346 => x"000000",
   23347 => x"000000",
   23348 => x"000000",
   23349 => x"00057f",
   23350 => x"ffffff",
   23351 => x"ffffff",
   23352 => x"ffffff",
   23353 => x"ffffd5",
   23354 => x"000015",
   23355 => x"aaaaaa",
   23356 => x"aaaa95",
   23357 => x"000000",
   23358 => x"015fff",
   23359 => x"ffffff",
   23360 => x"ffffff",
   23361 => x"ffffff",
   23362 => x"fffff5",
   23363 => x"c30c30",
   23364 => x"c30c30",
   23365 => x"c30c30",
   23366 => x"c30c30",
   23367 => x"c30c30",
   23368 => x"c30c30",
   23369 => x"c30c30",
   23370 => x"c30c30",
   23371 => x"c30c30",
   23372 => x"c30c30",
   23373 => x"c30c30",
   23374 => x"857df3",
   23375 => x"cf3cf3",
   23376 => x"cf3cf3",
   23377 => x"cf3cf3",
   23378 => x"cf3cf3",
   23379 => x"cf3cf3",
   23380 => x"cf3cf3",
   23381 => x"cf3cf3",
   23382 => x"cf3cf3",
   23383 => x"cf3cf3",
   23384 => x"cf3aae",
   23385 => x"ffffff",
   23386 => x"ffffff",
   23387 => x"ffffff",
   23388 => x"ffffff",
   23389 => x"ffffff",
   23390 => x"ffffff",
   23391 => x"ffffff",
   23392 => x"ffffff",
   23393 => x"ffffff",
   23394 => x"ffffff",
   23395 => x"ffffff",
   23396 => x"ffffff",
   23397 => x"ffffff",
   23398 => x"ffffff",
   23399 => x"ffffff",
   23400 => x"ffffff",
   23401 => x"ffffff",
   23402 => x"ffffff",
   23403 => x"ffffee",
   23404 => x"38f3cf",
   23405 => x"3cf3cf",
   23406 => x"3cf3cf",
   23407 => x"3cf3cf",
   23408 => x"3cf3cf",
   23409 => x"3cf3cf",
   23410 => x"3cf3cf",
   23411 => x"3cf3cf",
   23412 => x"3cf3cf",
   23413 => x"3cf3cf",
   23414 => x"3cd30c",
   23415 => x"30c30c",
   23416 => x"30c30c",
   23417 => x"30c30c",
   23418 => x"30c30c",
   23419 => x"30c30c",
   23420 => x"30c30c",
   23421 => x"30c30c",
   23422 => x"30c30c",
   23423 => x"30c30c",
   23424 => x"30c30c",
   23425 => x"30c32e",
   23426 => x"ffffff",
   23427 => x"ffffff",
   23428 => x"ffffff",
   23429 => x"ffffff",
   23430 => x"ffffff",
   23431 => x"ffffff",
   23432 => x"ffffff",
   23433 => x"ffffff",
   23434 => x"ffffff",
   23435 => x"a95abf",
   23436 => x"ffffff",
   23437 => x"ffffff",
   23438 => x"ffffff",
   23439 => x"ffffff",
   23440 => x"ffffff",
   23441 => x"fffeb0",
   23442 => x"c30c30",
   23443 => x"c30c30",
   23444 => x"c30c30",
   23445 => x"c30c30",
   23446 => x"c30c30",
   23447 => x"c30c30",
   23448 => x"c30c30",
   23449 => x"c30c30",
   23450 => x"c30c30",
   23451 => x"c30c30",
   23452 => x"c30c30",
   23453 => x"820820",
   23454 => x"820820",
   23455 => x"820820",
   23456 => x"820820",
   23457 => x"820820",
   23458 => x"820820",
   23459 => x"820820",
   23460 => x"820820",
   23461 => x"820820",
   23462 => x"820820",
   23463 => x"820820",
   23464 => x"820820",
   23465 => x"820820",
   23466 => x"820820",
   23467 => x"820820",
   23468 => x"820820",
   23469 => x"820820",
   23470 => x"820820",
   23471 => x"820820",
   23472 => x"820820",
   23473 => x"820820",
   23474 => x"820820",
   23475 => x"820410",
   23476 => x"410410",
   23477 => x"410410",
   23478 => x"410410",
   23479 => x"410410",
   23480 => x"410410",
   23481 => x"410410",
   23482 => x"410410",
   23483 => x"410410",
   23484 => x"410410",
   23485 => x"410410",
   23486 => x"410410",
   23487 => x"410410",
   23488 => x"410410",
   23489 => x"410410",
   23490 => x"410410",
   23491 => x"410410",
   23492 => x"410410",
   23493 => x"410410",
   23494 => x"410410",
   23495 => x"410410",
   23496 => x"410410",
   23497 => x"410410",
   23498 => x"410000",
   23499 => x"000000",
   23500 => x"000000",
   23501 => x"000000",
   23502 => x"000000",
   23503 => x"000000",
   23504 => x"000000",
   23505 => x"000000",
   23506 => x"000000",
   23507 => x"000000",
   23508 => x"000000",
   23509 => x"00057f",
   23510 => x"ffffff",
   23511 => x"ffffff",
   23512 => x"ffffff",
   23513 => x"ffffd5",
   23514 => x"00002a",
   23515 => x"ffffff",
   23516 => x"ffffff",
   23517 => x"a95000",
   23518 => x"000abf",
   23519 => x"ffffff",
   23520 => x"ffffff",
   23521 => x"ffffff",
   23522 => x"fffffa",
   23523 => x"c30c30",
   23524 => x"c30c30",
   23525 => x"c30c30",
   23526 => x"c30c30",
   23527 => x"c30c30",
   23528 => x"c30c30",
   23529 => x"c30c30",
   23530 => x"c30c30",
   23531 => x"c30c30",
   23532 => x"c30c30",
   23533 => x"c30c30",
   23534 => x"4a7cf3",
   23535 => x"cf3cf3",
   23536 => x"cf3cf3",
   23537 => x"cf3cf3",
   23538 => x"cf3cf3",
   23539 => x"cf3cf3",
   23540 => x"cf3cf3",
   23541 => x"cf3cf3",
   23542 => x"cf3cf3",
   23543 => x"cf3cf3",
   23544 => x"cf39ea",
   23545 => x"ffffff",
   23546 => x"ffffff",
   23547 => x"ffffff",
   23548 => x"ffffff",
   23549 => x"ffffff",
   23550 => x"ffffff",
   23551 => x"ffffff",
   23552 => x"ffffff",
   23553 => x"ffffff",
   23554 => x"ffffff",
   23555 => x"ffffff",
   23556 => x"ffffff",
   23557 => x"ffffff",
   23558 => x"ffffff",
   23559 => x"ffffff",
   23560 => x"ffffff",
   23561 => x"ffffff",
   23562 => x"ffffff",
   23563 => x"fffb9e",
   23564 => x"3cf3cf",
   23565 => x"3cf3cf",
   23566 => x"3cf3cf",
   23567 => x"3cf3cf",
   23568 => x"3cf3cf",
   23569 => x"3cf3cf",
   23570 => x"3cf3cf",
   23571 => x"3cf3cf",
   23572 => x"3cf3cf",
   23573 => x"3cf3cf",
   23574 => x"3ce30c",
   23575 => x"30c30c",
   23576 => x"30c30c",
   23577 => x"30c30c",
   23578 => x"30c30c",
   23579 => x"30c30c",
   23580 => x"30c30c",
   23581 => x"30c30c",
   23582 => x"30c30c",
   23583 => x"30c30c",
   23584 => x"30c30c",
   23585 => x"30c77f",
   23586 => x"ffffff",
   23587 => x"ffffff",
   23588 => x"ffffff",
   23589 => x"ffffff",
   23590 => x"ffffff",
   23591 => x"ffffff",
   23592 => x"ffffff",
   23593 => x"ffffff",
   23594 => x"ffffea",
   23595 => x"56afff",
   23596 => x"ffffff",
   23597 => x"ffffff",
   23598 => x"ffffff",
   23599 => x"ffffff",
   23600 => x"ffffff",
   23601 => x"fffeb0",
   23602 => x"c30c30",
   23603 => x"c30c30",
   23604 => x"c30c30",
   23605 => x"c30c30",
   23606 => x"c30c30",
   23607 => x"c30c30",
   23608 => x"c30c30",
   23609 => x"c30c30",
   23610 => x"c30c30",
   23611 => x"c30c30",
   23612 => x"c30c30",
   23613 => x"820820",
   23614 => x"820820",
   23615 => x"820820",
   23616 => x"820820",
   23617 => x"820820",
   23618 => x"820820",
   23619 => x"820820",
   23620 => x"820820",
   23621 => x"820820",
   23622 => x"820820",
   23623 => x"820820",
   23624 => x"820820",
   23625 => x"820820",
   23626 => x"820820",
   23627 => x"820820",
   23628 => x"820820",
   23629 => x"820820",
   23630 => x"820820",
   23631 => x"820820",
   23632 => x"820820",
   23633 => x"820820",
   23634 => x"820820",
   23635 => x"820410",
   23636 => x"410410",
   23637 => x"410410",
   23638 => x"410410",
   23639 => x"410410",
   23640 => x"410410",
   23641 => x"410410",
   23642 => x"410410",
   23643 => x"410410",
   23644 => x"410410",
   23645 => x"410410",
   23646 => x"410410",
   23647 => x"410410",
   23648 => x"410410",
   23649 => x"410410",
   23650 => x"410410",
   23651 => x"410410",
   23652 => x"410410",
   23653 => x"410410",
   23654 => x"410410",
   23655 => x"410410",
   23656 => x"410410",
   23657 => x"410410",
   23658 => x"410000",
   23659 => x"000000",
   23660 => x"000000",
   23661 => x"000000",
   23662 => x"000000",
   23663 => x"000000",
   23664 => x"000000",
   23665 => x"000000",
   23666 => x"000000",
   23667 => x"000000",
   23668 => x"000000",
   23669 => x"00057f",
   23670 => x"ffffff",
   23671 => x"ffffff",
   23672 => x"ffffff",
   23673 => x"ffffd5",
   23674 => x"00002a",
   23675 => x"ffffff",
   23676 => x"ffffff",
   23677 => x"fea000",
   23678 => x"00057f",
   23679 => x"ffffff",
   23680 => x"ffffff",
   23681 => x"ffffff",
   23682 => x"ffffff",
   23683 => x"d70c30",
   23684 => x"c30c30",
   23685 => x"c30c30",
   23686 => x"c30c30",
   23687 => x"c30c30",
   23688 => x"c30c30",
   23689 => x"c30c30",
   23690 => x"c30c30",
   23691 => x"c30c30",
   23692 => x"c30c30",
   23693 => x"c30c21",
   23694 => x"9f7cf3",
   23695 => x"cf3cf3",
   23696 => x"cf3cf3",
   23697 => x"cf3cf3",
   23698 => x"cf3cf3",
   23699 => x"cf3cf3",
   23700 => x"cf3cf3",
   23701 => x"cf3cf3",
   23702 => x"cf3cf3",
   23703 => x"cf3cf3",
   23704 => x"cf3ceb",
   23705 => x"bbffff",
   23706 => x"ffffff",
   23707 => x"ffffff",
   23708 => x"ffffff",
   23709 => x"ffffff",
   23710 => x"ffffff",
   23711 => x"ffffff",
   23712 => x"ffffff",
   23713 => x"ffffff",
   23714 => x"ffffff",
   23715 => x"ffffff",
   23716 => x"ffffff",
   23717 => x"ffffff",
   23718 => x"ffffff",
   23719 => x"ffffff",
   23720 => x"ffffff",
   23721 => x"ffffff",
   23722 => x"ffffff",
   23723 => x"fff78e",
   23724 => x"3cf3cf",
   23725 => x"3cf3cf",
   23726 => x"3cf3cf",
   23727 => x"3cf3cf",
   23728 => x"3cf3cf",
   23729 => x"3cf3cf",
   23730 => x"3cf3cf",
   23731 => x"3cf3cf",
   23732 => x"3cf3cf",
   23733 => x"3cf3cf",
   23734 => x"3cf34c",
   23735 => x"30c30c",
   23736 => x"30c30c",
   23737 => x"30c30c",
   23738 => x"30c30c",
   23739 => x"30c30c",
   23740 => x"30c30c",
   23741 => x"30c30c",
   23742 => x"30c30c",
   23743 => x"30c30c",
   23744 => x"30c30c",
   23745 => x"30cbbf",
   23746 => x"ffffff",
   23747 => x"ffffff",
   23748 => x"ffffff",
   23749 => x"ffffff",
   23750 => x"ffffff",
   23751 => x"ffffff",
   23752 => x"ffffff",
   23753 => x"ffffff",
   23754 => x"fffa95",
   23755 => x"abffff",
   23756 => x"ffffff",
   23757 => x"ffffff",
   23758 => x"ffffff",
   23759 => x"ffffff",
   23760 => x"ffffff",
   23761 => x"fffeb0",
   23762 => x"c30c30",
   23763 => x"c30c30",
   23764 => x"c30c30",
   23765 => x"c30c30",
   23766 => x"c30c30",
   23767 => x"c30c30",
   23768 => x"c30c30",
   23769 => x"c30c30",
   23770 => x"c30c30",
   23771 => x"c30c30",
   23772 => x"c30c30",
   23773 => x"820820",
   23774 => x"820820",
   23775 => x"820820",
   23776 => x"820820",
   23777 => x"820820",
   23778 => x"820820",
   23779 => x"820820",
   23780 => x"820820",
   23781 => x"820820",
   23782 => x"820820",
   23783 => x"820820",
   23784 => x"820820",
   23785 => x"820820",
   23786 => x"820820",
   23787 => x"820820",
   23788 => x"820820",
   23789 => x"820820",
   23790 => x"820820",
   23791 => x"820820",
   23792 => x"820820",
   23793 => x"820820",
   23794 => x"820820",
   23795 => x"820410",
   23796 => x"410410",
   23797 => x"410410",
   23798 => x"410410",
   23799 => x"410410",
   23800 => x"410410",
   23801 => x"410410",
   23802 => x"410410",
   23803 => x"410410",
   23804 => x"410410",
   23805 => x"410410",
   23806 => x"410410",
   23807 => x"410410",
   23808 => x"410410",
   23809 => x"410410",
   23810 => x"410410",
   23811 => x"410410",
   23812 => x"410410",
   23813 => x"410410",
   23814 => x"410410",
   23815 => x"410410",
   23816 => x"410410",
   23817 => x"410410",
   23818 => x"410000",
   23819 => x"000000",
   23820 => x"000000",
   23821 => x"000000",
   23822 => x"000000",
   23823 => x"000000",
   23824 => x"000000",
   23825 => x"000000",
   23826 => x"000000",
   23827 => x"000000",
   23828 => x"000000",
   23829 => x"00057f",
   23830 => x"ffffff",
   23831 => x"ffffff",
   23832 => x"ffffff",
   23833 => x"ffffd5",
   23834 => x"00002a",
   23835 => x"ffffff",
   23836 => x"ffffff",
   23837 => x"fff540",
   23838 => x"00057f",
   23839 => x"ffffff",
   23840 => x"ffffff",
   23841 => x"ffffff",
   23842 => x"ffffff",
   23843 => x"eb5c30",
   23844 => x"c30c30",
   23845 => x"c30c30",
   23846 => x"c30c30",
   23847 => x"c30c30",
   23848 => x"c30c30",
   23849 => x"c30c30",
   23850 => x"c30c30",
   23851 => x"c30c30",
   23852 => x"c30c30",
   23853 => x"c30c16",
   23854 => x"df3cf3",
   23855 => x"cf3cf3",
   23856 => x"cf3cf3",
   23857 => x"cf3cf3",
   23858 => x"cf3cf3",
   23859 => x"cf3cf3",
   23860 => x"cf3cf3",
   23861 => x"cf3cf3",
   23862 => x"cf3cf3",
   23863 => x"cf3cf3",
   23864 => x"cf3cf7",
   23865 => x"abffff",
   23866 => x"ffffff",
   23867 => x"ffffff",
   23868 => x"ffffff",
   23869 => x"ffffff",
   23870 => x"ffffff",
   23871 => x"ffffff",
   23872 => x"ffffff",
   23873 => x"ffffff",
   23874 => x"ffffff",
   23875 => x"ffffff",
   23876 => x"ffffff",
   23877 => x"ffffff",
   23878 => x"ffffff",
   23879 => x"ffffff",
   23880 => x"ffffff",
   23881 => x"ffffff",
   23882 => x"ffffff",
   23883 => x"fee78f",
   23884 => x"3cf3cf",
   23885 => x"3cf3cf",
   23886 => x"3cf3cf",
   23887 => x"3cf3cf",
   23888 => x"3cf3cf",
   23889 => x"3cf3cf",
   23890 => x"3cf3cf",
   23891 => x"3cf3cf",
   23892 => x"3cf3cf",
   23893 => x"3cf3cf",
   23894 => x"3cf38c",
   23895 => x"30c30c",
   23896 => x"30c30c",
   23897 => x"30c30c",
   23898 => x"30c30c",
   23899 => x"30c30c",
   23900 => x"30c30c",
   23901 => x"30c30c",
   23902 => x"30c30c",
   23903 => x"30c30c",
   23904 => x"30c30c",
   23905 => x"31dfff",
   23906 => x"ffffff",
   23907 => x"ffffff",
   23908 => x"ffffff",
   23909 => x"ffffff",
   23910 => x"ffffff",
   23911 => x"ffffff",
   23912 => x"ffffff",
   23913 => x"ffffff",
   23914 => x"fea56a",
   23915 => x"ffffff",
   23916 => x"ffffff",
   23917 => x"ffffff",
   23918 => x"ffffff",
   23919 => x"ffffff",
   23920 => x"ffffff",
   23921 => x"fffeb0",
   23922 => x"c30c30",
   23923 => x"c30c30",
   23924 => x"c30c30",
   23925 => x"c30c30",
   23926 => x"c30c30",
   23927 => x"c30c30",
   23928 => x"c30c30",
   23929 => x"c30c30",
   23930 => x"c30c30",
   23931 => x"c30c30",
   23932 => x"c30c30",
   23933 => x"820820",
   23934 => x"820820",
   23935 => x"820820",
   23936 => x"820820",
   23937 => x"820820",
   23938 => x"820820",
   23939 => x"820820",
   23940 => x"820820",
   23941 => x"820820",
   23942 => x"820820",
   23943 => x"820820",
   23944 => x"820820",
   23945 => x"820820",
   23946 => x"820820",
   23947 => x"820820",
   23948 => x"820820",
   23949 => x"820820",
   23950 => x"820820",
   23951 => x"820820",
   23952 => x"820820",
   23953 => x"820820",
   23954 => x"820820",
   23955 => x"820410",
   23956 => x"410410",
   23957 => x"410410",
   23958 => x"410410",
   23959 => x"410410",
   23960 => x"410410",
   23961 => x"410410",
   23962 => x"410410",
   23963 => x"410410",
   23964 => x"410410",
   23965 => x"410410",
   23966 => x"410410",
   23967 => x"410410",
   23968 => x"410410",
   23969 => x"410410",
   23970 => x"410410",
   23971 => x"410410",
   23972 => x"410410",
   23973 => x"410410",
   23974 => x"410410",
   23975 => x"410410",
   23976 => x"410410",
   23977 => x"410410",
   23978 => x"410000",
   23979 => x"000000",
   23980 => x"000000",
   23981 => x"000000",
   23982 => x"000000",
   23983 => x"000000",
   23984 => x"000000",
   23985 => x"000000",
   23986 => x"000000",
   23987 => x"000000",
   23988 => x"000000",
   23989 => x"00057f",
   23990 => x"ffffff",
   23991 => x"ffffff",
   23992 => x"ffffff",
   23993 => x"ffffd5",
   23994 => x"00002a",
   23995 => x"ffffff",
   23996 => x"ffffff",
   23997 => x"fff540",
   23998 => x"00057f",
   23999 => x"ffffff",
   24000 => x"ffffff",
   24001 => x"ffffff",
   24002 => x"ffffff",
   24003 => x"ffac30",
   24004 => x"c30c30",
   24005 => x"c30c30",
   24006 => x"c30c30",
   24007 => x"c30c30",
   24008 => x"c30c30",
   24009 => x"c30c30",
   24010 => x"c30c30",
   24011 => x"c30c30",
   24012 => x"c30c30",
   24013 => x"c3086b",
   24014 => x"cf3cf3",
   24015 => x"cf3cf3",
   24016 => x"cf3cf3",
   24017 => x"cf3cf3",
   24018 => x"cf3cf3",
   24019 => x"cf3cf3",
   24020 => x"cf3cf3",
   24021 => x"cf3cf3",
   24022 => x"cf3cf3",
   24023 => x"cf3cf3",
   24024 => x"cf3cf3",
   24025 => x"9eefff",
   24026 => x"ffffff",
   24027 => x"ffffff",
   24028 => x"ffffff",
   24029 => x"ffffff",
   24030 => x"ffffff",
   24031 => x"ffffff",
   24032 => x"ffffff",
   24033 => x"ffffff",
   24034 => x"ffffff",
   24035 => x"ffffff",
   24036 => x"ffffff",
   24037 => x"ffffff",
   24038 => x"ffffff",
   24039 => x"ffffff",
   24040 => x"ffffff",
   24041 => x"ffffff",
   24042 => x"ffffff",
   24043 => x"fde38f",
   24044 => x"3cf3cf",
   24045 => x"3cf3cf",
   24046 => x"3cf3cf",
   24047 => x"3cf3cf",
   24048 => x"3cf3cf",
   24049 => x"3cf3cf",
   24050 => x"3cf3cf",
   24051 => x"3cf3cf",
   24052 => x"3cf3cf",
   24053 => x"3cf3cf",
   24054 => x"3cf3cd",
   24055 => x"30c30c",
   24056 => x"30c30c",
   24057 => x"30c30c",
   24058 => x"30c30c",
   24059 => x"30c30c",
   24060 => x"30c30c",
   24061 => x"30c30c",
   24062 => x"30c30c",
   24063 => x"30c30c",
   24064 => x"30c30c",
   24065 => x"76efff",
   24066 => x"ffffff",
   24067 => x"ffffff",
   24068 => x"ffffff",
   24069 => x"ffffff",
   24070 => x"ffffff",
   24071 => x"ffffff",
   24072 => x"ffffff",
   24073 => x"ffffff",
   24074 => x"a95abf",
   24075 => x"ffffff",
   24076 => x"ffffff",
   24077 => x"ffffff",
   24078 => x"ffffff",
   24079 => x"ffffff",
   24080 => x"ffffff",
   24081 => x"fffeb0",
   24082 => x"c30c30",
   24083 => x"c30c30",
   24084 => x"c30c30",
   24085 => x"c30c30",
   24086 => x"c30c30",
   24087 => x"c30c30",
   24088 => x"c30c30",
   24089 => x"c30c30",
   24090 => x"c30c30",
   24091 => x"c30c30",
   24092 => x"c30c30",
   24093 => x"820820",
   24094 => x"820820",
   24095 => x"820820",
   24096 => x"820820",
   24097 => x"820820",
   24098 => x"820820",
   24099 => x"820820",
   24100 => x"820820",
   24101 => x"820820",
   24102 => x"820820",
   24103 => x"820820",
   24104 => x"820820",
   24105 => x"820820",
   24106 => x"820820",
   24107 => x"820820",
   24108 => x"820820",
   24109 => x"820820",
   24110 => x"820820",
   24111 => x"820820",
   24112 => x"820820",
   24113 => x"820820",
   24114 => x"820820",
   24115 => x"820410",
   24116 => x"410410",
   24117 => x"410410",
   24118 => x"410410",
   24119 => x"410410",
   24120 => x"410410",
   24121 => x"410410",
   24122 => x"410410",
   24123 => x"410410",
   24124 => x"410410",
   24125 => x"410410",
   24126 => x"410410",
   24127 => x"410410",
   24128 => x"410410",
   24129 => x"410410",
   24130 => x"410410",
   24131 => x"410410",
   24132 => x"410410",
   24133 => x"410410",
   24134 => x"410410",
   24135 => x"410410",
   24136 => x"410410",
   24137 => x"410410",
   24138 => x"410000",
   24139 => x"000000",
   24140 => x"000000",
   24141 => x"000000",
   24142 => x"000000",
   24143 => x"000000",
   24144 => x"000000",
   24145 => x"000000",
   24146 => x"000000",
   24147 => x"000000",
   24148 => x"000000",
   24149 => x"00057f",
   24150 => x"ffffff",
   24151 => x"ffffff",
   24152 => x"ffffff",
   24153 => x"ffffd5",
   24154 => x"00002a",
   24155 => x"ffffff",
   24156 => x"ffffff",
   24157 => x"fffa80",
   24158 => x"00057f",
   24159 => x"ffffff",
   24160 => x"ffffff",
   24161 => x"ffffff",
   24162 => x"ffffff",
   24163 => x"ffad70",
   24164 => x"c30c30",
   24165 => x"c30c30",
   24166 => x"c30c30",
   24167 => x"c30c30",
   24168 => x"c30c30",
   24169 => x"c30c30",
   24170 => x"c30c30",
   24171 => x"c30c30",
   24172 => x"c30c30",
   24173 => x"c305b7",
   24174 => x"cf3cf3",
   24175 => x"cf3cf3",
   24176 => x"cf3cf3",
   24177 => x"cf3cf3",
   24178 => x"cf3cf3",
   24179 => x"cf3cf3",
   24180 => x"cf3cf3",
   24181 => x"cf3cf3",
   24182 => x"cf3cf3",
   24183 => x"cf3cf3",
   24184 => x"cf3cf3",
   24185 => x"ceabbf",
   24186 => x"ffffff",
   24187 => x"ffffff",
   24188 => x"ffffff",
   24189 => x"ffffff",
   24190 => x"ffffff",
   24191 => x"ffffff",
   24192 => x"ffffff",
   24193 => x"ffffff",
   24194 => x"ffffff",
   24195 => x"ffffff",
   24196 => x"ffffff",
   24197 => x"ffffff",
   24198 => x"ffffff",
   24199 => x"ffffff",
   24200 => x"ffffff",
   24201 => x"ffffff",
   24202 => x"ffffff",
   24203 => x"b9e3cf",
   24204 => x"3cf3cf",
   24205 => x"3cf3cf",
   24206 => x"3cf3cf",
   24207 => x"3cf3cf",
   24208 => x"3cf3cf",
   24209 => x"3cf3cf",
   24210 => x"3cf3cf",
   24211 => x"3cf3cf",
   24212 => x"3cf3cf",
   24213 => x"3cf3cf",
   24214 => x"3cf3ce",
   24215 => x"30c30c",
   24216 => x"30c30c",
   24217 => x"30c30c",
   24218 => x"30c30c",
   24219 => x"30c30c",
   24220 => x"30c30c",
   24221 => x"30c30c",
   24222 => x"30c30c",
   24223 => x"30c30c",
   24224 => x"30c30c",
   24225 => x"77ffff",
   24226 => x"ffffff",
   24227 => x"ffffff",
   24228 => x"ffffff",
   24229 => x"ffffff",
   24230 => x"ffffff",
   24231 => x"ffffff",
   24232 => x"ffffff",
   24233 => x"ffffea",
   24234 => x"56afff",
   24235 => x"ffffff",
   24236 => x"ffffff",
   24237 => x"ffffff",
   24238 => x"ffffff",
   24239 => x"ffffff",
   24240 => x"ffffff",
   24241 => x"fffeb0",
   24242 => x"c30c30",
   24243 => x"c30c30",
   24244 => x"c30c30",
   24245 => x"c30c30",
   24246 => x"c30c30",
   24247 => x"c30c30",
   24248 => x"c30c30",
   24249 => x"c30c30",
   24250 => x"c30c30",
   24251 => x"c30c30",
   24252 => x"c30c30",
   24253 => x"820820",
   24254 => x"820820",
   24255 => x"820820",
   24256 => x"820820",
   24257 => x"820820",
   24258 => x"820820",
   24259 => x"820820",
   24260 => x"820820",
   24261 => x"820820",
   24262 => x"820820",
   24263 => x"820820",
   24264 => x"820820",
   24265 => x"820820",
   24266 => x"820820",
   24267 => x"820820",
   24268 => x"820820",
   24269 => x"820820",
   24270 => x"820820",
   24271 => x"820820",
   24272 => x"820820",
   24273 => x"820820",
   24274 => x"820820",
   24275 => x"820410",
   24276 => x"410410",
   24277 => x"410410",
   24278 => x"410410",
   24279 => x"410410",
   24280 => x"410410",
   24281 => x"410410",
   24282 => x"410410",
   24283 => x"410410",
   24284 => x"410410",
   24285 => x"410410",
   24286 => x"410410",
   24287 => x"410410",
   24288 => x"410410",
   24289 => x"410410",
   24290 => x"410410",
   24291 => x"410410",
   24292 => x"410410",
   24293 => x"410410",
   24294 => x"410410",
   24295 => x"410410",
   24296 => x"410410",
   24297 => x"410410",
   24298 => x"410000",
   24299 => x"000000",
   24300 => x"000000",
   24301 => x"000000",
   24302 => x"000000",
   24303 => x"000000",
   24304 => x"000000",
   24305 => x"000000",
   24306 => x"000000",
   24307 => x"000000",
   24308 => x"000000",
   24309 => x"00057f",
   24310 => x"ffffff",
   24311 => x"ffffff",
   24312 => x"ffffff",
   24313 => x"ffffd5",
   24314 => x"00002a",
   24315 => x"ffffff",
   24316 => x"ffffff",
   24317 => x"fff540",
   24318 => x"00057f",
   24319 => x"ffffff",
   24320 => x"ffffff",
   24321 => x"ffffff",
   24322 => x"ffffff",
   24323 => x"fffeb0",
   24324 => x"c30c30",
   24325 => x"c30c30",
   24326 => x"c30c30",
   24327 => x"c30c30",
   24328 => x"c30c30",
   24329 => x"c30c30",
   24330 => x"c30c30",
   24331 => x"c30c30",
   24332 => x"c30c30",
   24333 => x"c219f3",
   24334 => x"cf3cf3",
   24335 => x"cf3cf3",
   24336 => x"cf3cf3",
   24337 => x"cf3cf3",
   24338 => x"cf3cf3",
   24339 => x"cf3cf3",
   24340 => x"cf3cf3",
   24341 => x"cf3cf3",
   24342 => x"cf3cf3",
   24343 => x"cf3cf3",
   24344 => x"cf3cf3",
   24345 => x"cf7bbf",
   24346 => x"ffffff",
   24347 => x"ffffff",
   24348 => x"ffffff",
   24349 => x"ffffff",
   24350 => x"ffffff",
   24351 => x"ffffff",
   24352 => x"ffffff",
   24353 => x"ffffff",
   24354 => x"ffffff",
   24355 => x"ffffff",
   24356 => x"ffffff",
   24357 => x"ffffff",
   24358 => x"ffffff",
   24359 => x"ffffff",
   24360 => x"ffffff",
   24361 => x"ffffff",
   24362 => x"ffffff",
   24363 => x"78e3cf",
   24364 => x"3cf3cf",
   24365 => x"3cf3cf",
   24366 => x"3cf3cf",
   24367 => x"3cf3cf",
   24368 => x"3cf3cf",
   24369 => x"3cf3cf",
   24370 => x"3cf3cf",
   24371 => x"3cf3cf",
   24372 => x"3cf3cf",
   24373 => x"3cf3cf",
   24374 => x"3cf3cf",
   24375 => x"34c30c",
   24376 => x"30c30c",
   24377 => x"30c30c",
   24378 => x"30c30c",
   24379 => x"30c30c",
   24380 => x"30c30c",
   24381 => x"30c30c",
   24382 => x"30c30c",
   24383 => x"30c30c",
   24384 => x"30c31d",
   24385 => x"ffffff",
   24386 => x"ffffff",
   24387 => x"ffffff",
   24388 => x"ffffff",
   24389 => x"ffffff",
   24390 => x"ffffff",
   24391 => x"ffffff",
   24392 => x"ffffff",
   24393 => x"fffa95",
   24394 => x"abffff",
   24395 => x"ffffff",
   24396 => x"ffffff",
   24397 => x"ffffff",
   24398 => x"ffffff",
   24399 => x"ffffff",
   24400 => x"ffffff",
   24401 => x"fffeb0",
   24402 => x"c30c30",
   24403 => x"c30c30",
   24404 => x"c30c30",
   24405 => x"c30c30",
   24406 => x"c30c30",
   24407 => x"c30c30",
   24408 => x"c30c30",
   24409 => x"c30c30",
   24410 => x"c30c30",
   24411 => x"c30c30",
   24412 => x"c30c30",
   24413 => x"820820",
   24414 => x"820820",
   24415 => x"820820",
   24416 => x"820820",
   24417 => x"820820",
   24418 => x"820820",
   24419 => x"820820",
   24420 => x"820820",
   24421 => x"820820",
   24422 => x"820820",
   24423 => x"820820",
   24424 => x"820820",
   24425 => x"820820",
   24426 => x"820820",
   24427 => x"820820",
   24428 => x"820820",
   24429 => x"820820",
   24430 => x"820820",
   24431 => x"820820",
   24432 => x"820820",
   24433 => x"820820",
   24434 => x"820820",
   24435 => x"820410",
   24436 => x"410410",
   24437 => x"410410",
   24438 => x"410410",
   24439 => x"410410",
   24440 => x"410410",
   24441 => x"410410",
   24442 => x"410410",
   24443 => x"410410",
   24444 => x"410410",
   24445 => x"410410",
   24446 => x"410410",
   24447 => x"410410",
   24448 => x"410410",
   24449 => x"410410",
   24450 => x"410410",
   24451 => x"410410",
   24452 => x"410410",
   24453 => x"410410",
   24454 => x"410410",
   24455 => x"410410",
   24456 => x"410410",
   24457 => x"410410",
   24458 => x"410000",
   24459 => x"000000",
   24460 => x"000000",
   24461 => x"000000",
   24462 => x"000000",
   24463 => x"000000",
   24464 => x"000000",
   24465 => x"000000",
   24466 => x"000000",
   24467 => x"000000",
   24468 => x"000000",
   24469 => x"00057f",
   24470 => x"ffffff",
   24471 => x"ffffff",
   24472 => x"ffffff",
   24473 => x"ffffd5",
   24474 => x"00002a",
   24475 => x"ffffff",
   24476 => x"ffffff",
   24477 => x"fea540",
   24478 => x"00057f",
   24479 => x"ffffff",
   24480 => x"ffffff",
   24481 => x"ffffff",
   24482 => x"ffffff",
   24483 => x"fffff5",
   24484 => x"c30c30",
   24485 => x"c30c30",
   24486 => x"c30c30",
   24487 => x"c30c30",
   24488 => x"c30c30",
   24489 => x"c30c30",
   24490 => x"c30c30",
   24491 => x"c30c30",
   24492 => x"c30c30",
   24493 => x"c12df3",
   24494 => x"cf3cf3",
   24495 => x"cf3cf3",
   24496 => x"cf3cf3",
   24497 => x"cf3cf3",
   24498 => x"cf3cf3",
   24499 => x"cf3cf3",
   24500 => x"cf3cf3",
   24501 => x"cf3cf3",
   24502 => x"cf3cf3",
   24503 => x"cf3cf3",
   24504 => x"cf3cf3",
   24505 => x"cf3aee",
   24506 => x"ffffff",
   24507 => x"ffffff",
   24508 => x"ffffff",
   24509 => x"ffffff",
   24510 => x"ffffff",
   24511 => x"ffffff",
   24512 => x"ffffff",
   24513 => x"ffffff",
   24514 => x"ffffff",
   24515 => x"ffffff",
   24516 => x"ffffff",
   24517 => x"ffffff",
   24518 => x"ffffff",
   24519 => x"ffffff",
   24520 => x"ffffff",
   24521 => x"ffffff",
   24522 => x"ffffee",
   24523 => x"38f3cf",
   24524 => x"3cf3cf",
   24525 => x"3cf3cf",
   24526 => x"3cf3cf",
   24527 => x"3cf3cf",
   24528 => x"3cf3cf",
   24529 => x"3cf3cf",
   24530 => x"3cf3cf",
   24531 => x"3cf3cf",
   24532 => x"3cf3cf",
   24533 => x"3cf3cf",
   24534 => x"3cf3cf",
   24535 => x"38c30c",
   24536 => x"30c30c",
   24537 => x"30c30c",
   24538 => x"30c30c",
   24539 => x"30c30c",
   24540 => x"30c30c",
   24541 => x"30c30c",
   24542 => x"30c30c",
   24543 => x"30c30c",
   24544 => x"30c32e",
   24545 => x"ffffff",
   24546 => x"ffffff",
   24547 => x"ffffff",
   24548 => x"ffffff",
   24549 => x"ffffff",
   24550 => x"ffffff",
   24551 => x"ffffff",
   24552 => x"ffffff",
   24553 => x"fea56a",
   24554 => x"ffffff",
   24555 => x"ffffff",
   24556 => x"ffffff",
   24557 => x"ffffff",
   24558 => x"ffffff",
   24559 => x"ffffff",
   24560 => x"ffffff",
   24561 => x"fffeb0",
   24562 => x"c30c30",
   24563 => x"c30c30",
   24564 => x"c30c30",
   24565 => x"c30c30",
   24566 => x"c30c30",
   24567 => x"c30c30",
   24568 => x"c30c30",
   24569 => x"c30c30",
   24570 => x"c30c30",
   24571 => x"c30c30",
   24572 => x"c30c30",
   24573 => x"820820",
   24574 => x"820820",
   24575 => x"820820",
   24576 => x"820820",
   24577 => x"820820",
   24578 => x"820820",
   24579 => x"820820",
   24580 => x"820820",
   24581 => x"820820",
   24582 => x"820820",
   24583 => x"820820",
   24584 => x"820820",
   24585 => x"820820",
   24586 => x"820820",
   24587 => x"820820",
   24588 => x"820820",
   24589 => x"820820",
   24590 => x"820820",
   24591 => x"820820",
   24592 => x"820820",
   24593 => x"820820",
   24594 => x"820820",
   24595 => x"820410",
   24596 => x"410410",
   24597 => x"410410",
   24598 => x"410410",
   24599 => x"410410",
   24600 => x"410410",
   24601 => x"410410",
   24602 => x"410410",
   24603 => x"410410",
   24604 => x"410410",
   24605 => x"410410",
   24606 => x"410410",
   24607 => x"410410",
   24608 => x"410410",
   24609 => x"410410",
   24610 => x"410410",
   24611 => x"410410",
   24612 => x"410410",
   24613 => x"410410",
   24614 => x"410410",
   24615 => x"410410",
   24616 => x"410410",
   24617 => x"410410",
   24618 => x"410000",
   24619 => x"000000",
   24620 => x"000000",
   24621 => x"000000",
   24622 => x"000000",
   24623 => x"000000",
   24624 => x"000000",
   24625 => x"000000",
   24626 => x"000000",
   24627 => x"000000",
   24628 => x"000000",
   24629 => x"00057f",
   24630 => x"ffffff",
   24631 => x"ffffff",
   24632 => x"ffffff",
   24633 => x"ffffd5",
   24634 => x"00002a",
   24635 => x"ffffff",
   24636 => x"ffffff",
   24637 => x"fea000",
   24638 => x"000abf",
   24639 => x"ffffff",
   24640 => x"ffffff",
   24641 => x"ffffff",
   24642 => x"ffffff",
   24643 => x"fffffa",
   24644 => x"d70c30",
   24645 => x"c30c30",
   24646 => x"c30c30",
   24647 => x"c30c30",
   24648 => x"c30c30",
   24649 => x"c30c30",
   24650 => x"c30c30",
   24651 => x"c30c30",
   24652 => x"c30c30",
   24653 => x"867cf3",
   24654 => x"cf3cf3",
   24655 => x"cf3cf3",
   24656 => x"cf3cf3",
   24657 => x"cf3cf3",
   24658 => x"cf3cf3",
   24659 => x"cf3cf3",
   24660 => x"cf3cf3",
   24661 => x"cf3cf3",
   24662 => x"cf3cf3",
   24663 => x"cf3cf3",
   24664 => x"cf3cf3",
   24665 => x"cf3dda",
   24666 => x"ffffff",
   24667 => x"ffffff",
   24668 => x"ffffff",
   24669 => x"ffffff",
   24670 => x"ffffff",
   24671 => x"ffffff",
   24672 => x"ffffff",
   24673 => x"ffffff",
   24674 => x"ffffff",
   24675 => x"ffffff",
   24676 => x"ffffff",
   24677 => x"ffffff",
   24678 => x"ffffff",
   24679 => x"ffffff",
   24680 => x"ffffff",
   24681 => x"ffffff",
   24682 => x"fffb9e",
   24683 => x"3cf3cf",
   24684 => x"3cf3cf",
   24685 => x"3cf3cf",
   24686 => x"3cf3cf",
   24687 => x"3cf3cf",
   24688 => x"3cf3cf",
   24689 => x"3cf3cf",
   24690 => x"3cf3cf",
   24691 => x"3cf3cf",
   24692 => x"3cf3cf",
   24693 => x"3cf3cf",
   24694 => x"3cf3cf",
   24695 => x"3cd30c",
   24696 => x"30c30c",
   24697 => x"30c30c",
   24698 => x"30c30c",
   24699 => x"30c30c",
   24700 => x"30c30c",
   24701 => x"30c30c",
   24702 => x"30c30c",
   24703 => x"30c30c",
   24704 => x"30c77f",
   24705 => x"ffffff",
   24706 => x"ffffff",
   24707 => x"ffffff",
   24708 => x"ffffff",
   24709 => x"ffffff",
   24710 => x"ffffff",
   24711 => x"ffffff",
   24712 => x"ffffff",
   24713 => x"a95abf",
   24714 => x"ffffff",
   24715 => x"ffffff",
   24716 => x"ffffff",
   24717 => x"ffffff",
   24718 => x"ffffff",
   24719 => x"ffffff",
   24720 => x"ffffff",
   24721 => x"fffeb0",
   24722 => x"c30c30",
   24723 => x"c30c30",
   24724 => x"c30c30",
   24725 => x"c30c30",
   24726 => x"c30c30",
   24727 => x"c30c30",
   24728 => x"c30c30",
   24729 => x"c30c30",
   24730 => x"c30c30",
   24731 => x"c30c30",
   24732 => x"c30c30",
   24733 => x"820820",
   24734 => x"820820",
   24735 => x"820820",
   24736 => x"820820",
   24737 => x"820820",
   24738 => x"820820",
   24739 => x"820820",
   24740 => x"820820",
   24741 => x"820820",
   24742 => x"820820",
   24743 => x"820820",
   24744 => x"820820",
   24745 => x"820820",
   24746 => x"820820",
   24747 => x"820820",
   24748 => x"820820",
   24749 => x"820820",
   24750 => x"820820",
   24751 => x"820820",
   24752 => x"820820",
   24753 => x"820820",
   24754 => x"820820",
   24755 => x"820410",
   24756 => x"410410",
   24757 => x"410410",
   24758 => x"410410",
   24759 => x"410410",
   24760 => x"410410",
   24761 => x"410410",
   24762 => x"410410",
   24763 => x"410410",
   24764 => x"410410",
   24765 => x"410410",
   24766 => x"410410",
   24767 => x"410410",
   24768 => x"410410",
   24769 => x"410410",
   24770 => x"410410",
   24771 => x"410410",
   24772 => x"410410",
   24773 => x"410410",
   24774 => x"410410",
   24775 => x"410410",
   24776 => x"410410",
   24777 => x"410410",
   24778 => x"410000",
   24779 => x"000000",
   24780 => x"000000",
   24781 => x"000000",
   24782 => x"000000",
   24783 => x"000000",
   24784 => x"000000",
   24785 => x"000000",
   24786 => x"000000",
   24787 => x"000000",
   24788 => x"000000",
   24789 => x"00057f",
   24790 => x"ffffff",
   24791 => x"ffffff",
   24792 => x"ffffff",
   24793 => x"ffffd5",
   24794 => x"00002a",
   24795 => x"ffffff",
   24796 => x"ffffff",
   24797 => x"a95000",
   24798 => x"015fff",
   24799 => x"ffffff",
   24800 => x"ffffff",
   24801 => x"ffffff",
   24802 => x"ffffff",
   24803 => x"ffffff",
   24804 => x"eb0c30",
   24805 => x"c30c30",
   24806 => x"c30c30",
   24807 => x"c30c30",
   24808 => x"c30c30",
   24809 => x"c30c30",
   24810 => x"c30c30",
   24811 => x"c30c30",
   24812 => x"c30c30",
   24813 => x"4b7cf3",
   24814 => x"cf3cf3",
   24815 => x"cf3cf3",
   24816 => x"cf3cf3",
   24817 => x"cf3cf3",
   24818 => x"cf3cf3",
   24819 => x"cf3cf3",
   24820 => x"cf3cf3",
   24821 => x"cf3cf3",
   24822 => x"cf3cf3",
   24823 => x"cf3cf3",
   24824 => x"cf3cf3",
   24825 => x"cf3ce7",
   24826 => x"bbffff",
   24827 => x"ffffff",
   24828 => x"ffffff",
   24829 => x"ffffff",
   24830 => x"ffffff",
   24831 => x"ffffff",
   24832 => x"ffffff",
   24833 => x"ffffff",
   24834 => x"ffffff",
   24835 => x"ffffff",
   24836 => x"ffffff",
   24837 => x"ffffff",
   24838 => x"ffffff",
   24839 => x"ffffff",
   24840 => x"ffffff",
   24841 => x"ffffff",
   24842 => x"fff78e",
   24843 => x"3cf3cf",
   24844 => x"3cf3cf",
   24845 => x"3cf3cf",
   24846 => x"3cf3cf",
   24847 => x"3cf3cf",
   24848 => x"3cf3cf",
   24849 => x"3cf3cf",
   24850 => x"3cf3cf",
   24851 => x"3cf3cf",
   24852 => x"3cf3cf",
   24853 => x"3cf3cf",
   24854 => x"3cf3cf",
   24855 => x"3ce30c",
   24856 => x"30c30c",
   24857 => x"30c30c",
   24858 => x"30c30c",
   24859 => x"30c30c",
   24860 => x"30c30c",
   24861 => x"30c30c",
   24862 => x"30c30c",
   24863 => x"30c30c",
   24864 => x"31dbbf",
   24865 => x"ffffff",
   24866 => x"ffffff",
   24867 => x"ffffff",
   24868 => x"ffffff",
   24869 => x"ffffff",
   24870 => x"ffffff",
   24871 => x"ffffff",
   24872 => x"ffffea",
   24873 => x"56afff",
   24874 => x"ffffff",
   24875 => x"ffffff",
   24876 => x"ffffff",
   24877 => x"ffffff",
   24878 => x"ffffff",
   24879 => x"ffffff",
   24880 => x"ffffff",
   24881 => x"fffeb0",
   24882 => x"c30c30",
   24883 => x"c30c30",
   24884 => x"c30c30",
   24885 => x"c30c30",
   24886 => x"c30c30",
   24887 => x"c30c30",
   24888 => x"c30c30",
   24889 => x"c30c30",
   24890 => x"c30c30",
   24891 => x"c30c30",
   24892 => x"c30c30",
   24893 => x"820820",
   24894 => x"820820",
   24895 => x"820820",
   24896 => x"820820",
   24897 => x"820820",
   24898 => x"820820",
   24899 => x"820820",
   24900 => x"820820",
   24901 => x"820820",
   24902 => x"820820",
   24903 => x"820820",
   24904 => x"820820",
   24905 => x"820820",
   24906 => x"820820",
   24907 => x"820820",
   24908 => x"820820",
   24909 => x"820820",
   24910 => x"820820",
   24911 => x"820820",
   24912 => x"820820",
   24913 => x"820820",
   24914 => x"820820",
   24915 => x"820410",
   24916 => x"410410",
   24917 => x"410410",
   24918 => x"410410",
   24919 => x"410410",
   24920 => x"410410",
   24921 => x"410410",
   24922 => x"410410",
   24923 => x"410410",
   24924 => x"410410",
   24925 => x"410410",
   24926 => x"410410",
   24927 => x"410410",
   24928 => x"410410",
   24929 => x"410410",
   24930 => x"410410",
   24931 => x"410410",
   24932 => x"410410",
   24933 => x"410410",
   24934 => x"410410",
   24935 => x"410410",
   24936 => x"410410",
   24937 => x"410410",
   24938 => x"410000",
   24939 => x"000000",
   24940 => x"000000",
   24941 => x"000000",
   24942 => x"000000",
   24943 => x"000000",
   24944 => x"000000",
   24945 => x"000000",
   24946 => x"000000",
   24947 => x"000000",
   24948 => x"000000",
   24949 => x"00057f",
   24950 => x"ffffff",
   24951 => x"ffffff",
   24952 => x"ffffff",
   24953 => x"ffffd5",
   24954 => x"00002a",
   24955 => x"abffff",
   24956 => x"aaaa95",
   24957 => x"000000",
   24958 => x"56afff",
   24959 => x"ffffff",
   24960 => x"ffffff",
   24961 => x"ffffff",
   24962 => x"ffffff",
   24963 => x"ffffff",
   24964 => x"ff5c30",
   24965 => x"c30c30",
   24966 => x"c30c30",
   24967 => x"c30c30",
   24968 => x"c30c30",
   24969 => x"c30c30",
   24970 => x"c30c30",
   24971 => x"c30c30",
   24972 => x"c30c30",
   24973 => x"5f7cf3",
   24974 => x"cf3cf3",
   24975 => x"cf3cf3",
   24976 => x"cf3cf3",
   24977 => x"cf3cf3",
   24978 => x"cf3cf3",
   24979 => x"cf3cf3",
   24980 => x"cf3cf3",
   24981 => x"cf3cf3",
   24982 => x"cf3cf3",
   24983 => x"cf3cf3",
   24984 => x"cf3cf3",
   24985 => x"cf3cf3",
   24986 => x"aaefff",
   24987 => x"ffffff",
   24988 => x"ffffff",
   24989 => x"ffffff",
   24990 => x"ffffff",
   24991 => x"ffffff",
   24992 => x"ffffff",
   24993 => x"ffffff",
   24994 => x"ffffff",
   24995 => x"ffffff",
   24996 => x"ffffff",
   24997 => x"ffffff",
   24998 => x"ffffff",
   24999 => x"ffffff",
   25000 => x"ffffff",
   25001 => x"ffffff",
   25002 => x"fdd38f",
   25003 => x"3cf3cf",
   25004 => x"3cf3cf",
   25005 => x"3cf3cf",
   25006 => x"3cf3cf",
   25007 => x"3cf3cf",
   25008 => x"3cf3cf",
   25009 => x"3cf3cf",
   25010 => x"3cf3cf",
   25011 => x"3cf3cf",
   25012 => x"3cf3cf",
   25013 => x"3cf3cf",
   25014 => x"3cf3cf",
   25015 => x"3ce34c",
   25016 => x"30c30c",
   25017 => x"30c30c",
   25018 => x"30c30c",
   25019 => x"30c30c",
   25020 => x"30c30c",
   25021 => x"30c30c",
   25022 => x"30c30c",
   25023 => x"30c30c",
   25024 => x"32efff",
   25025 => x"ffffff",
   25026 => x"ffffff",
   25027 => x"ffffff",
   25028 => x"ffffff",
   25029 => x"ffffff",
   25030 => x"ffffff",
   25031 => x"ffffff",
   25032 => x"fffa95",
   25033 => x"abffff",
   25034 => x"ffffff",
   25035 => x"ffffff",
   25036 => x"ffffff",
   25037 => x"ffffff",
   25038 => x"ffffff",
   25039 => x"ffffff",
   25040 => x"ffffff",
   25041 => x"fffeb0",
   25042 => x"c30c30",
   25043 => x"c30c30",
   25044 => x"c30c30",
   25045 => x"c30c30",
   25046 => x"c30c30",
   25047 => x"c30c30",
   25048 => x"c30c30",
   25049 => x"c30c30",
   25050 => x"c30c30",
   25051 => x"c30c30",
   25052 => x"c30c30",
   25053 => x"820820",
   25054 => x"820820",
   25055 => x"820820",
   25056 => x"820820",
   25057 => x"820820",
   25058 => x"820820",
   25059 => x"820820",
   25060 => x"820820",
   25061 => x"820820",
   25062 => x"820820",
   25063 => x"820820",
   25064 => x"820820",
   25065 => x"820820",
   25066 => x"820820",
   25067 => x"820820",
   25068 => x"820820",
   25069 => x"820820",
   25070 => x"820820",
   25071 => x"820820",
   25072 => x"820820",
   25073 => x"820820",
   25074 => x"820820",
   25075 => x"820410",
   25076 => x"410410",
   25077 => x"410410",
   25078 => x"410410",
   25079 => x"410410",
   25080 => x"410410",
   25081 => x"410410",
   25082 => x"410410",
   25083 => x"410410",
   25084 => x"410410",
   25085 => x"410410",
   25086 => x"410410",
   25087 => x"410410",
   25088 => x"410410",
   25089 => x"410410",
   25090 => x"410410",
   25091 => x"410410",
   25092 => x"410410",
   25093 => x"410410",
   25094 => x"410410",
   25095 => x"410410",
   25096 => x"410410",
   25097 => x"410410",
   25098 => x"410000",
   25099 => x"000000",
   25100 => x"000000",
   25101 => x"000000",
   25102 => x"000000",
   25103 => x"000000",
   25104 => x"000000",
   25105 => x"000000",
   25106 => x"000000",
   25107 => x"000000",
   25108 => x"000000",
   25109 => x"00057f",
   25110 => x"ffffff",
   25111 => x"ffffff",
   25112 => x"ffffff",
   25113 => x"ffffd5",
   25114 => x"000000",
   25115 => x"000000",
   25116 => x"000000",
   25117 => x"000015",
   25118 => x"abffff",
   25119 => x"ffffff",
   25120 => x"ffffff",
   25121 => x"ffffff",
   25122 => x"ffffff",
   25123 => x"ffffff",
   25124 => x"ffad70",
   25125 => x"c30c30",
   25126 => x"c30c30",
   25127 => x"c30c30",
   25128 => x"c30c30",
   25129 => x"c30c30",
   25130 => x"c30c30",
   25131 => x"c30c30",
   25132 => x"c30c21",
   25133 => x"9f3cf3",
   25134 => x"cf3cf3",
   25135 => x"cf3cf3",
   25136 => x"cf3cf3",
   25137 => x"cf3cf3",
   25138 => x"cf3cf3",
   25139 => x"cf3cf3",
   25140 => x"cf3cf3",
   25141 => x"cf3cf3",
   25142 => x"cf3cf3",
   25143 => x"cf3cf3",
   25144 => x"cf3cf3",
   25145 => x"cf3cf3",
   25146 => x"ddafff",
   25147 => x"ffffff",
   25148 => x"ffffff",
   25149 => x"ffffff",
   25150 => x"ffffff",
   25151 => x"ffffff",
   25152 => x"ffffff",
   25153 => x"ffffff",
   25154 => x"ffffff",
   25155 => x"ffffff",
   25156 => x"ffffff",
   25157 => x"ffffff",
   25158 => x"ffffff",
   25159 => x"ffffff",
   25160 => x"ffffff",
   25161 => x"ffffff",
   25162 => x"b8e3cf",
   25163 => x"3cf3cf",
   25164 => x"3cf3cf",
   25165 => x"3cf3cf",
   25166 => x"3cf3cf",
   25167 => x"3cf3cf",
   25168 => x"3cf3cf",
   25169 => x"3cf3cf",
   25170 => x"3cf3cf",
   25171 => x"3cf3cf",
   25172 => x"3cf3cf",
   25173 => x"3cf3cf",
   25174 => x"3cf3cf",
   25175 => x"3cf34c",
   25176 => x"30c30c",
   25177 => x"30c30c",
   25178 => x"30c30c",
   25179 => x"30c30c",
   25180 => x"30c30c",
   25181 => x"30c30c",
   25182 => x"30c30c",
   25183 => x"30c30c",
   25184 => x"77ffff",
   25185 => x"ffffff",
   25186 => x"ffffff",
   25187 => x"ffffff",
   25188 => x"ffffff",
   25189 => x"ffffff",
   25190 => x"ffffff",
   25191 => x"ffffff",
   25192 => x"fea56a",
   25193 => x"ffffff",
   25194 => x"ffffff",
   25195 => x"ffffff",
   25196 => x"ffffff",
   25197 => x"ffffff",
   25198 => x"ffffff",
   25199 => x"ffffff",
   25200 => x"ffffff",
   25201 => x"fffeb0",
   25202 => x"c30c30",
   25203 => x"c30c30",
   25204 => x"c30c30",
   25205 => x"c30c30",
   25206 => x"c30c30",
   25207 => x"c30c30",
   25208 => x"c30c30",
   25209 => x"c30c30",
   25210 => x"c30c30",
   25211 => x"c30c30",
   25212 => x"c30c30",
   25213 => x"820820",
   25214 => x"820820",
   25215 => x"820820",
   25216 => x"820820",
   25217 => x"820820",
   25218 => x"820820",
   25219 => x"820820",
   25220 => x"820820",
   25221 => x"820820",
   25222 => x"820820",
   25223 => x"820820",
   25224 => x"820820",
   25225 => x"820820",
   25226 => x"820820",
   25227 => x"820820",
   25228 => x"820820",
   25229 => x"820820",
   25230 => x"820820",
   25231 => x"820820",
   25232 => x"820820",
   25233 => x"820820",
   25234 => x"820820",
   25235 => x"820410",
   25236 => x"410410",
   25237 => x"410410",
   25238 => x"410410",
   25239 => x"410410",
   25240 => x"410410",
   25241 => x"410410",
   25242 => x"410410",
   25243 => x"410410",
   25244 => x"410410",
   25245 => x"410410",
   25246 => x"410410",
   25247 => x"410410",
   25248 => x"410410",
   25249 => x"410410",
   25250 => x"410410",
   25251 => x"410410",
   25252 => x"410410",
   25253 => x"410410",
   25254 => x"410410",
   25255 => x"410410",
   25256 => x"410410",
   25257 => x"410410",
   25258 => x"410000",
   25259 => x"000000",
   25260 => x"000000",
   25261 => x"000000",
   25262 => x"000000",
   25263 => x"000000",
   25264 => x"000000",
   25265 => x"000000",
   25266 => x"000000",
   25267 => x"000000",
   25268 => x"000000",
   25269 => x"00057f",
   25270 => x"ffffff",
   25271 => x"ffffff",
   25272 => x"ffffff",
   25273 => x"ffffd5",
   25274 => x"000000",
   25275 => x"000000",
   25276 => x"000000",
   25277 => x"00057f",
   25278 => x"ffffff",
   25279 => x"ffffff",
   25280 => x"ffffff",
   25281 => x"ffffff",
   25282 => x"ffffff",
   25283 => x"ffffff",
   25284 => x"fffeb0",
   25285 => x"c30c30",
   25286 => x"c30c30",
   25287 => x"c30c30",
   25288 => x"c30c30",
   25289 => x"c30c30",
   25290 => x"c30c30",
   25291 => x"c30c30",
   25292 => x"c30c12",
   25293 => x"df3cf3",
   25294 => x"cf3cf3",
   25295 => x"cf3cf3",
   25296 => x"cf3cf3",
   25297 => x"cf3cf3",
   25298 => x"cf3cf3",
   25299 => x"cf3cf3",
   25300 => x"cf3cf3",
   25301 => x"cf3cf3",
   25302 => x"cf3cf3",
   25303 => x"cf3cf3",
   25304 => x"cf3cf3",
   25305 => x"cf3cf3",
   25306 => x"cf77bf",
   25307 => x"ffffff",
   25308 => x"ffffff",
   25309 => x"ffffff",
   25310 => x"ffffff",
   25311 => x"ffffff",
   25312 => x"ffffff",
   25313 => x"ffffff",
   25314 => x"ffffff",
   25315 => x"ffffff",
   25316 => x"ffffff",
   25317 => x"ffffff",
   25318 => x"ffffff",
   25319 => x"ffffff",
   25320 => x"ffffff",
   25321 => x"ffffee",
   25322 => x"74e3cf",
   25323 => x"3cf3cf",
   25324 => x"3cf3cf",
   25325 => x"3cf3cf",
   25326 => x"3cf3cf",
   25327 => x"3cf3cf",
   25328 => x"3cf3cf",
   25329 => x"3cf3cf",
   25330 => x"3cf3cf",
   25331 => x"3cf3cf",
   25332 => x"3cf3cf",
   25333 => x"3cf3cf",
   25334 => x"3cf3cf",
   25335 => x"3cf38d",
   25336 => x"30c30c",
   25337 => x"30c30c",
   25338 => x"30c30c",
   25339 => x"30c30c",
   25340 => x"30c30c",
   25341 => x"30c30c",
   25342 => x"30c30c",
   25343 => x"30c31d",
   25344 => x"bbffff",
   25345 => x"ffffff",
   25346 => x"ffffff",
   25347 => x"ffffff",
   25348 => x"ffffff",
   25349 => x"ffffff",
   25350 => x"ffffff",
   25351 => x"ffffff",
   25352 => x"a95abf",
   25353 => x"ffffff",
   25354 => x"ffffff",
   25355 => x"ffffff",
   25356 => x"ffffff",
   25357 => x"ffffff",
   25358 => x"ffffff",
   25359 => x"ffffff",
   25360 => x"ffffff",
   25361 => x"fffeb0",
   25362 => x"c30c30",
   25363 => x"c30c30",
   25364 => x"c30c30",
   25365 => x"c30c30",
   25366 => x"c30c30",
   25367 => x"c30c30",
   25368 => x"c30c30",
   25369 => x"c30c30",
   25370 => x"c30c30",
   25371 => x"c30c30",
   25372 => x"c30c30",
   25373 => x"820820",
   25374 => x"820820",
   25375 => x"820820",
   25376 => x"820820",
   25377 => x"820820",
   25378 => x"820820",
   25379 => x"820820",
   25380 => x"820820",
   25381 => x"820820",
   25382 => x"820820",
   25383 => x"820820",
   25384 => x"820820",
   25385 => x"820820",
   25386 => x"820820",
   25387 => x"820820",
   25388 => x"820820",
   25389 => x"820820",
   25390 => x"820820",
   25391 => x"820820",
   25392 => x"820820",
   25393 => x"820820",
   25394 => x"820820",
   25395 => x"820410",
   25396 => x"410410",
   25397 => x"410410",
   25398 => x"410410",
   25399 => x"410410",
   25400 => x"410410",
   25401 => x"410410",
   25402 => x"410410",
   25403 => x"410410",
   25404 => x"410410",
   25405 => x"410410",
   25406 => x"410410",
   25407 => x"410410",
   25408 => x"410410",
   25409 => x"410410",
   25410 => x"410410",
   25411 => x"410410",
   25412 => x"410410",
   25413 => x"410410",
   25414 => x"410410",
   25415 => x"410410",
   25416 => x"410410",
   25417 => x"410410",
   25418 => x"410000",
   25419 => x"000000",
   25420 => x"000000",
   25421 => x"000000",
   25422 => x"000000",
   25423 => x"000000",
   25424 => x"000000",
   25425 => x"000000",
   25426 => x"000000",
   25427 => x"000000",
   25428 => x"000000",
   25429 => x"00057f",
   25430 => x"ffffff",
   25431 => x"ffffff",
   25432 => x"ffffff",
   25433 => x"ffffd5",
   25434 => x"000000",
   25435 => x"000000",
   25436 => x"000000",
   25437 => x"00056a",
   25438 => x"ffffff",
   25439 => x"ffffff",
   25440 => x"ffffff",
   25441 => x"ffffff",
   25442 => x"ffffff",
   25443 => x"ffffff",
   25444 => x"fffffa",
   25445 => x"c30c30",
   25446 => x"c30c30",
   25447 => x"c30c30",
   25448 => x"c30c30",
   25449 => x"c30c30",
   25450 => x"c30c30",
   25451 => x"c30c30",
   25452 => x"c30867",
   25453 => x"cf3cf3",
   25454 => x"cf3cf3",
   25455 => x"cf3cf3",
   25456 => x"cf3cf3",
   25457 => x"cf3cf3",
   25458 => x"cf3cf3",
   25459 => x"cf3cf3",
   25460 => x"cf3cf3",
   25461 => x"cf3cf3",
   25462 => x"cf3cf3",
   25463 => x"cf3cf3",
   25464 => x"cf3cf3",
   25465 => x"cf3cf3",
   25466 => x"cf3aee",
   25467 => x"ffffff",
   25468 => x"ffffff",
   25469 => x"ffffff",
   25470 => x"ffffff",
   25471 => x"ffffff",
   25472 => x"ffffff",
   25473 => x"ffffff",
   25474 => x"ffffff",
   25475 => x"ffffff",
   25476 => x"ffffff",
   25477 => x"ffffff",
   25478 => x"ffffff",
   25479 => x"ffffff",
   25480 => x"ffffff",
   25481 => x"ffffdd",
   25482 => x"38f3cf",
   25483 => x"3cf3cf",
   25484 => x"3cf3cf",
   25485 => x"3cf3cf",
   25486 => x"3cf3cf",
   25487 => x"3cf3cf",
   25488 => x"3cf3cf",
   25489 => x"3cf3cf",
   25490 => x"3cf3cf",
   25491 => x"3cf3cf",
   25492 => x"3cf3cf",
   25493 => x"3cf3cf",
   25494 => x"3cf3cf",
   25495 => x"3cf3cd",
   25496 => x"30c30c",
   25497 => x"30c30c",
   25498 => x"30c30c",
   25499 => x"30c30c",
   25500 => x"30c30c",
   25501 => x"30c30c",
   25502 => x"30c30c",
   25503 => x"30c76e",
   25504 => x"ffffff",
   25505 => x"ffffff",
   25506 => x"ffffff",
   25507 => x"ffffff",
   25508 => x"ffffff",
   25509 => x"ffffff",
   25510 => x"ffffff",
   25511 => x"ffffea",
   25512 => x"56afff",
   25513 => x"ffffff",
   25514 => x"ffffff",
   25515 => x"ffffff",
   25516 => x"ffffff",
   25517 => x"ffffff",
   25518 => x"ffffff",
   25519 => x"ffffff",
   25520 => x"ffffff",
   25521 => x"fffeb0",
   25522 => x"c30c30",
   25523 => x"c30c30",
   25524 => x"c30c30",
   25525 => x"c30c30",
   25526 => x"c30c30",
   25527 => x"c30c30",
   25528 => x"c30c30",
   25529 => x"c30c30",
   25530 => x"c30c30",
   25531 => x"c30c30",
   25532 => x"c30c30",
   25533 => x"820820",
   25534 => x"820820",
   25535 => x"820820",
   25536 => x"820820",
   25537 => x"820820",
   25538 => x"820820",
   25539 => x"820820",
   25540 => x"820820",
   25541 => x"820820",
   25542 => x"820820",
   25543 => x"820820",
   25544 => x"820820",
   25545 => x"820820",
   25546 => x"820820",
   25547 => x"820820",
   25548 => x"820820",
   25549 => x"820820",
   25550 => x"820820",
   25551 => x"820820",
   25552 => x"820820",
   25553 => x"820820",
   25554 => x"820820",
   25555 => x"820410",
   25556 => x"410410",
   25557 => x"410410",
   25558 => x"410410",
   25559 => x"410410",
   25560 => x"410410",
   25561 => x"410410",
   25562 => x"410410",
   25563 => x"410410",
   25564 => x"410410",
   25565 => x"410410",
   25566 => x"410410",
   25567 => x"410410",
   25568 => x"410410",
   25569 => x"410410",
   25570 => x"410410",
   25571 => x"410410",
   25572 => x"410410",
   25573 => x"410410",
   25574 => x"410410",
   25575 => x"410410",
   25576 => x"410410",
   25577 => x"410410",
   25578 => x"410000",
   25579 => x"000000",
   25580 => x"000000",
   25581 => x"000000",
   25582 => x"000000",
   25583 => x"000000",
   25584 => x"000000",
   25585 => x"000000",
   25586 => x"000000",
   25587 => x"000000",
   25588 => x"000000",
   25589 => x"00057f",
   25590 => x"ffffff",
   25591 => x"ffffff",
   25592 => x"ffffff",
   25593 => x"ffffd5",
   25594 => x"00002a",
   25595 => x"aaaaaa",
   25596 => x"aaa540",
   25597 => x"000015",
   25598 => x"abffff",
   25599 => x"ffffff",
   25600 => x"ffffff",
   25601 => x"ffffff",
   25602 => x"ffffff",
   25603 => x"ffffff",
   25604 => x"ffffff",
   25605 => x"d70c30",
   25606 => x"c30c30",
   25607 => x"c30c30",
   25608 => x"c30c30",
   25609 => x"c30c30",
   25610 => x"c30c30",
   25611 => x"c30c30",
   25612 => x"c308b7",
   25613 => x"cf3cf3",
   25614 => x"cf3cf3",
   25615 => x"cf3cf3",
   25616 => x"cf3cf3",
   25617 => x"cf3cf3",
   25618 => x"cf3cf3",
   25619 => x"cf3cf3",
   25620 => x"cf3cf3",
   25621 => x"cf3cf3",
   25622 => x"cf3cf3",
   25623 => x"cf3cf3",
   25624 => x"cf3cf3",
   25625 => x"cf3cf3",
   25626 => x"cf3cea",
   25627 => x"bfffff",
   25628 => x"ffffff",
   25629 => x"ffffff",
   25630 => x"ffffff",
   25631 => x"ffffff",
   25632 => x"ffffff",
   25633 => x"ffffff",
   25634 => x"ffffff",
   25635 => x"ffffff",
   25636 => x"ffffff",
   25637 => x"ffffff",
   25638 => x"ffffff",
   25639 => x"ffffff",
   25640 => x"ffffff",
   25641 => x"fff78e",
   25642 => x"3cf3cf",
   25643 => x"3cf3cf",
   25644 => x"3cf3cf",
   25645 => x"3cf3cf",
   25646 => x"3cf3cf",
   25647 => x"3cf3cf",
   25648 => x"3cf3cf",
   25649 => x"3cf3cf",
   25650 => x"3cf3cf",
   25651 => x"3cf3cf",
   25652 => x"3cf3cf",
   25653 => x"3cf3cf",
   25654 => x"3cf3cf",
   25655 => x"3cf3ce",
   25656 => x"30c30c",
   25657 => x"30c30c",
   25658 => x"30c30c",
   25659 => x"30c30c",
   25660 => x"30c30c",
   25661 => x"30c30c",
   25662 => x"30c30c",
   25663 => x"30cbbf",
   25664 => x"ffffff",
   25665 => x"ffffff",
   25666 => x"ffffff",
   25667 => x"ffffff",
   25668 => x"ffffff",
   25669 => x"ffffff",
   25670 => x"ffffff",
   25671 => x"fffa95",
   25672 => x"abffff",
   25673 => x"ffffff",
   25674 => x"ffffff",
   25675 => x"ffffff",
   25676 => x"ffffff",
   25677 => x"ffffff",
   25678 => x"ffffff",
   25679 => x"ffffff",
   25680 => x"ffffff",
   25681 => x"fffeb0",
   25682 => x"c30c30",
   25683 => x"c30c30",
   25684 => x"c30c30",
   25685 => x"c30c30",
   25686 => x"c30c30",
   25687 => x"c30c30",
   25688 => x"c30c30",
   25689 => x"c30c30",
   25690 => x"c30c30",
   25691 => x"c30c30",
   25692 => x"c30c30",
   25693 => x"820820",
   25694 => x"820820",
   25695 => x"820820",
   25696 => x"820820",
   25697 => x"820820",
   25698 => x"820820",
   25699 => x"820820",
   25700 => x"820820",
   25701 => x"820820",
   25702 => x"820820",
   25703 => x"820820",
   25704 => x"820820",
   25705 => x"820820",
   25706 => x"820820",
   25707 => x"820820",
   25708 => x"820820",
   25709 => x"820820",
   25710 => x"820820",
   25711 => x"820820",
   25712 => x"820820",
   25713 => x"820820",
   25714 => x"820820",
   25715 => x"820410",
   25716 => x"410410",
   25717 => x"410410",
   25718 => x"410410",
   25719 => x"410410",
   25720 => x"410410",
   25721 => x"410410",
   25722 => x"410410",
   25723 => x"410410",
   25724 => x"410410",
   25725 => x"410410",
   25726 => x"410410",
   25727 => x"410410",
   25728 => x"410410",
   25729 => x"410410",
   25730 => x"410410",
   25731 => x"410410",
   25732 => x"410410",
   25733 => x"410410",
   25734 => x"410410",
   25735 => x"410410",
   25736 => x"410410",
   25737 => x"410410",
   25738 => x"410000",
   25739 => x"000000",
   25740 => x"000000",
   25741 => x"000000",
   25742 => x"000000",
   25743 => x"000000",
   25744 => x"000000",
   25745 => x"000000",
   25746 => x"000000",
   25747 => x"000000",
   25748 => x"000000",
   25749 => x"00057f",
   25750 => x"ffffff",
   25751 => x"ffffff",
   25752 => x"ffffff",
   25753 => x"ffffd5",
   25754 => x"00002a",
   25755 => x"ffffff",
   25756 => x"ffffea",
   25757 => x"540000",
   25758 => x"57ffff",
   25759 => x"ffffff",
   25760 => x"ffffff",
   25761 => x"ffffff",
   25762 => x"ffffff",
   25763 => x"ffffff",
   25764 => x"ffffff",
   25765 => x"eb5c30",
   25766 => x"c30c30",
   25767 => x"c30c30",
   25768 => x"c30c30",
   25769 => x"c30c30",
   25770 => x"c30c30",
   25771 => x"c30c30",
   25772 => x"c305f7",
   25773 => x"cf3cf3",
   25774 => x"cf3cf3",
   25775 => x"cf3cf3",
   25776 => x"cf3cf3",
   25777 => x"cf3cf3",
   25778 => x"cf3cf3",
   25779 => x"cf3cf3",
   25780 => x"cf3cf3",
   25781 => x"cf3cf3",
   25782 => x"cf3cf3",
   25783 => x"cf3cf3",
   25784 => x"cf3cf3",
   25785 => x"cf3cf3",
   25786 => x"cf3cf7",
   25787 => x"6bffff",
   25788 => x"ffffff",
   25789 => x"ffffff",
   25790 => x"ffffff",
   25791 => x"ffffff",
   25792 => x"ffffff",
   25793 => x"ffffff",
   25794 => x"ffffff",
   25795 => x"ffffff",
   25796 => x"ffffff",
   25797 => x"ffffff",
   25798 => x"ffffff",
   25799 => x"ffffff",
   25800 => x"ffffff",
   25801 => x"fee38f",
   25802 => x"3cf3cf",
   25803 => x"3cf3cf",
   25804 => x"3cf3cf",
   25805 => x"3cf3cf",
   25806 => x"3cf3cf",
   25807 => x"3cf3cf",
   25808 => x"3cf3cf",
   25809 => x"3cf3cf",
   25810 => x"3cf3cf",
   25811 => x"3cf3cf",
   25812 => x"3cf3cf",
   25813 => x"3cf3cf",
   25814 => x"3cf3cf",
   25815 => x"3cf3ce",
   25816 => x"34c30c",
   25817 => x"30c30c",
   25818 => x"30c30c",
   25819 => x"30c30c",
   25820 => x"30c30c",
   25821 => x"30c30c",
   25822 => x"30c30c",
   25823 => x"31dfff",
   25824 => x"ffffff",
   25825 => x"ffffff",
   25826 => x"ffffff",
   25827 => x"ffffff",
   25828 => x"ffffff",
   25829 => x"ffffff",
   25830 => x"ffffff",
   25831 => x"fea56a",
   25832 => x"ffffff",
   25833 => x"ffffff",
   25834 => x"ffffff",
   25835 => x"ffffff",
   25836 => x"ffffff",
   25837 => x"ffffff",
   25838 => x"ffffff",
   25839 => x"ffffff",
   25840 => x"ffffff",
   25841 => x"fffeb0",
   25842 => x"c30c30",
   25843 => x"c30c30",
   25844 => x"c30c30",
   25845 => x"c30c30",
   25846 => x"c30c30",
   25847 => x"c30c30",
   25848 => x"c30c30",
   25849 => x"c30c30",
   25850 => x"c30c30",
   25851 => x"c30c30",
   25852 => x"c30c30",
   25853 => x"820820",
   25854 => x"820820",
   25855 => x"820820",
   25856 => x"820820",
   25857 => x"820820",
   25858 => x"820820",
   25859 => x"820820",
   25860 => x"820820",
   25861 => x"820820",
   25862 => x"820820",
   25863 => x"820820",
   25864 => x"820820",
   25865 => x"820820",
   25866 => x"820820",
   25867 => x"820820",
   25868 => x"820820",
   25869 => x"820820",
   25870 => x"820820",
   25871 => x"820820",
   25872 => x"820820",
   25873 => x"820820",
   25874 => x"820820",
   25875 => x"820410",
   25876 => x"410410",
   25877 => x"410410",
   25878 => x"410410",
   25879 => x"410410",
   25880 => x"410410",
   25881 => x"410410",
   25882 => x"410410",
   25883 => x"410410",
   25884 => x"410410",
   25885 => x"410410",
   25886 => x"410410",
   25887 => x"410410",
   25888 => x"410410",
   25889 => x"410410",
   25890 => x"410410",
   25891 => x"410410",
   25892 => x"410410",
   25893 => x"410410",
   25894 => x"410410",
   25895 => x"410410",
   25896 => x"410410",
   25897 => x"410410",
   25898 => x"410000",
   25899 => x"000000",
   25900 => x"000000",
   25901 => x"000000",
   25902 => x"000000",
   25903 => x"000000",
   25904 => x"000000",
   25905 => x"000000",
   25906 => x"000000",
   25907 => x"000000",
   25908 => x"000000",
   25909 => x"00057f",
   25910 => x"ffffff",
   25911 => x"ffffff",
   25912 => x"ffffff",
   25913 => x"ffffd5",
   25914 => x"00002a",
   25915 => x"ffffff",
   25916 => x"ffffff",
   25917 => x"a95000",
   25918 => x"015fff",
   25919 => x"ffffff",
   25920 => x"ffffff",
   25921 => x"ffffff",
   25922 => x"ffffff",
   25923 => x"ffffff",
   25924 => x"ffffff",
   25925 => x"ffac30",
   25926 => x"c30c30",
   25927 => x"c30c30",
   25928 => x"c30c30",
   25929 => x"c30c30",
   25930 => x"c30c30",
   25931 => x"c30c30",
   25932 => x"c219f3",
   25933 => x"cf3cf3",
   25934 => x"cf3cf3",
   25935 => x"cf3cf3",
   25936 => x"cf3cf3",
   25937 => x"cf3cf3",
   25938 => x"cf3cf3",
   25939 => x"cf3cf3",
   25940 => x"cf3cf3",
   25941 => x"cf3cf3",
   25942 => x"cf3cf3",
   25943 => x"cf3cf3",
   25944 => x"cf3cf3",
   25945 => x"cf3cf3",
   25946 => x"cf3cf3",
   25947 => x"9defff",
   25948 => x"ffffff",
   25949 => x"ffffff",
   25950 => x"ffffff",
   25951 => x"ffffff",
   25952 => x"ffffff",
   25953 => x"ffffff",
   25954 => x"ffffff",
   25955 => x"ffffff",
   25956 => x"ffffff",
   25957 => x"ffffff",
   25958 => x"ffffff",
   25959 => x"ffffff",
   25960 => x"ffffff",
   25961 => x"b8d3cf",
   25962 => x"3cf3cf",
   25963 => x"3cf3cf",
   25964 => x"3cf3cf",
   25965 => x"3cf3cf",
   25966 => x"3cf3cf",
   25967 => x"3cf3cf",
   25968 => x"3cf3cf",
   25969 => x"3cf3cf",
   25970 => x"3cf3cf",
   25971 => x"3cf3cf",
   25972 => x"3cf3cf",
   25973 => x"3cf3cf",
   25974 => x"3cf3cf",
   25975 => x"3cf3cf",
   25976 => x"34c30c",
   25977 => x"30c30c",
   25978 => x"30c30c",
   25979 => x"30c30c",
   25980 => x"30c30c",
   25981 => x"30c30c",
   25982 => x"30c30c",
   25983 => x"76efff",
   25984 => x"ffffff",
   25985 => x"ffffff",
   25986 => x"ffffff",
   25987 => x"ffffff",
   25988 => x"ffffff",
   25989 => x"ffffff",
   25990 => x"ffffff",
   25991 => x"a95abf",
   25992 => x"ffffff",
   25993 => x"ffffff",
   25994 => x"ffffff",
   25995 => x"ffffff",
   25996 => x"ffffff",
   25997 => x"ffffff",
   25998 => x"ffffff",
   25999 => x"ffffff",
   26000 => x"ffffff",
   26001 => x"fffeb0",
   26002 => x"c30c30",
   26003 => x"c30c30",
   26004 => x"c30c30",
   26005 => x"c30c30",
   26006 => x"c30c30",
   26007 => x"c30c30",
   26008 => x"c30c30",
   26009 => x"c30c30",
   26010 => x"c30c30",
   26011 => x"c30c30",
   26012 => x"c30c30",
   26013 => x"820820",
   26014 => x"820820",
   26015 => x"820820",
   26016 => x"820820",
   26017 => x"820820",
   26018 => x"820820",
   26019 => x"820820",
   26020 => x"820820",
   26021 => x"820820",
   26022 => x"820820",
   26023 => x"820820",
   26024 => x"820820",
   26025 => x"820820",
   26026 => x"820820",
   26027 => x"820820",
   26028 => x"820820",
   26029 => x"820820",
   26030 => x"820820",
   26031 => x"820820",
   26032 => x"820820",
   26033 => x"820820",
   26034 => x"820820",
   26035 => x"820410",
   26036 => x"410410",
   26037 => x"410410",
   26038 => x"410410",
   26039 => x"410410",
   26040 => x"410410",
   26041 => x"410410",
   26042 => x"410410",
   26043 => x"410410",
   26044 => x"410410",
   26045 => x"410410",
   26046 => x"410410",
   26047 => x"410410",
   26048 => x"410410",
   26049 => x"410410",
   26050 => x"410410",
   26051 => x"410410",
   26052 => x"410410",
   26053 => x"410410",
   26054 => x"410410",
   26055 => x"410410",
   26056 => x"410410",
   26057 => x"410410",
   26058 => x"410000",
   26059 => x"000000",
   26060 => x"000000",
   26061 => x"000000",
   26062 => x"000000",
   26063 => x"000000",
   26064 => x"000000",
   26065 => x"000000",
   26066 => x"000000",
   26067 => x"000000",
   26068 => x"000000",
   26069 => x"00057f",
   26070 => x"ffffff",
   26071 => x"ffffff",
   26072 => x"ffffff",
   26073 => x"ffffd5",
   26074 => x"00002a",
   26075 => x"ffffff",
   26076 => x"ffffff",
   26077 => x"fea000",
   26078 => x"015abf",
   26079 => x"ffffff",
   26080 => x"ffffff",
   26081 => x"ffffff",
   26082 => x"ffffff",
   26083 => x"ffffff",
   26084 => x"ffffff",
   26085 => x"fffeb0",
   26086 => x"c30c30",
   26087 => x"c30c30",
   26088 => x"c30c30",
   26089 => x"c30c30",
   26090 => x"c30c30",
   26091 => x"c30c30",
   26092 => x"c22df3",
   26093 => x"cf3cf3",
   26094 => x"cf3cf3",
   26095 => x"cf3cf3",
   26096 => x"cf3cf3",
   26097 => x"cf3cf3",
   26098 => x"cf3cf3",
   26099 => x"cf3cf3",
   26100 => x"cf3cf3",
   26101 => x"cf3cf3",
   26102 => x"cf3cf3",
   26103 => x"cf3cf3",
   26104 => x"cf3cf3",
   26105 => x"cf3cf3",
   26106 => x"cf3cf3",
   26107 => x"ce7bbf",
   26108 => x"ffffff",
   26109 => x"ffffff",
   26110 => x"ffffff",
   26111 => x"ffffff",
   26112 => x"ffffff",
   26113 => x"ffffff",
   26114 => x"ffffff",
   26115 => x"ffffff",
   26116 => x"ffffff",
   26117 => x"ffffff",
   26118 => x"ffffff",
   26119 => x"ffffff",
   26120 => x"ffffee",
   26121 => x"74e3cf",
   26122 => x"3cf3cf",
   26123 => x"3cf3cf",
   26124 => x"3cf3cf",
   26125 => x"3cf3cf",
   26126 => x"3cf3cf",
   26127 => x"3cf3cf",
   26128 => x"3cf3cf",
   26129 => x"3cf3cf",
   26130 => x"3cf3cf",
   26131 => x"3cf3cf",
   26132 => x"3cf3cf",
   26133 => x"3cf3cf",
   26134 => x"3cf3cf",
   26135 => x"3cf3cf",
   26136 => x"38c30c",
   26137 => x"30c30c",
   26138 => x"30c30c",
   26139 => x"30c30c",
   26140 => x"30c30c",
   26141 => x"30c30c",
   26142 => x"30c31d",
   26143 => x"bbffff",
   26144 => x"ffffff",
   26145 => x"ffffff",
   26146 => x"ffffff",
   26147 => x"ffffff",
   26148 => x"ffffff",
   26149 => x"ffffff",
   26150 => x"ffffea",
   26151 => x"56afff",
   26152 => x"ffffff",
   26153 => x"ffffff",
   26154 => x"ffffff",
   26155 => x"ffffff",
   26156 => x"ffffff",
   26157 => x"ffffff",
   26158 => x"ffffff",
   26159 => x"ffffff",
   26160 => x"ffffff",
   26161 => x"fffeb0",
   26162 => x"c30c30",
   26163 => x"c30c30",
   26164 => x"c30c30",
   26165 => x"c30c30",
   26166 => x"c30c30",
   26167 => x"c30c30",
   26168 => x"c30c30",
   26169 => x"c30c30",
   26170 => x"c30c30",
   26171 => x"c30c30",
   26172 => x"c30c30",
   26173 => x"820820",
   26174 => x"820820",
   26175 => x"820820",
   26176 => x"820820",
   26177 => x"820820",
   26178 => x"820820",
   26179 => x"820820",
   26180 => x"820820",
   26181 => x"820820",
   26182 => x"820820",
   26183 => x"820820",
   26184 => x"820820",
   26185 => x"820820",
   26186 => x"820820",
   26187 => x"820820",
   26188 => x"820820",
   26189 => x"820820",
   26190 => x"820820",
   26191 => x"820820",
   26192 => x"820820",
   26193 => x"820820",
   26194 => x"820820",
   26195 => x"820410",
   26196 => x"410410",
   26197 => x"410410",
   26198 => x"410410",
   26199 => x"410410",
   26200 => x"410410",
   26201 => x"410410",
   26202 => x"410410",
   26203 => x"410410",
   26204 => x"410410",
   26205 => x"410410",
   26206 => x"410410",
   26207 => x"410410",
   26208 => x"410410",
   26209 => x"410410",
   26210 => x"410410",
   26211 => x"410410",
   26212 => x"410410",
   26213 => x"410410",
   26214 => x"410410",
   26215 => x"410410",
   26216 => x"410410",
   26217 => x"410410",
   26218 => x"410000",
   26219 => x"000000",
   26220 => x"000000",
   26221 => x"000000",
   26222 => x"000000",
   26223 => x"000000",
   26224 => x"000000",
   26225 => x"000000",
   26226 => x"000000",
   26227 => x"000000",
   26228 => x"000000",
   26229 => x"00057f",
   26230 => x"ffffff",
   26231 => x"ffffff",
   26232 => x"ffffff",
   26233 => x"ffffd5",
   26234 => x"00002a",
   26235 => x"ffffff",
   26236 => x"ffffff",
   26237 => x"fea540",
   26238 => x"00057f",
   26239 => x"ffffff",
   26240 => x"ffffff",
   26241 => x"ffffff",
   26242 => x"ffffff",
   26243 => x"ffffff",
   26244 => x"ffffff",
   26245 => x"fffff5",
   26246 => x"c30c30",
   26247 => x"c30c30",
   26248 => x"c30c30",
   26249 => x"c30c30",
   26250 => x"c30c30",
   26251 => x"c30c30",
   26252 => x"c17df3",
   26253 => x"cf3cf3",
   26254 => x"cf3cf3",
   26255 => x"cf3cf3",
   26256 => x"cf3cf3",
   26257 => x"cf3cf3",
   26258 => x"cf3cf3",
   26259 => x"cf3cf3",
   26260 => x"cf3cf3",
   26261 => x"cf3cf3",
   26262 => x"cf3cf3",
   26263 => x"cf3cf3",
   26264 => x"cf3cf3",
   26265 => x"cf3cf3",
   26266 => x"cf3cf3",
   26267 => x"cf3aae",
   26268 => x"ffffff",
   26269 => x"ffffff",
   26270 => x"ffffff",
   26271 => x"ffffff",
   26272 => x"ffffff",
   26273 => x"ffffff",
   26274 => x"ffffff",
   26275 => x"ffffff",
   26276 => x"ffffff",
   26277 => x"ffffff",
   26278 => x"ffffff",
   26279 => x"ffffff",
   26280 => x"fffb9d",
   26281 => x"38f3cf",
   26282 => x"3cf3cf",
   26283 => x"3cf3cf",
   26284 => x"3cf3cf",
   26285 => x"3cf3cf",
   26286 => x"3cf3cf",
   26287 => x"3cf3cf",
   26288 => x"3cf3cf",
   26289 => x"3cf3cf",
   26290 => x"3cf3cf",
   26291 => x"3cf3cf",
   26292 => x"3cf3cf",
   26293 => x"3cf3cf",
   26294 => x"3cf3cf",
   26295 => x"3cf3cf",
   26296 => x"38d30c",
   26297 => x"30c30c",
   26298 => x"30c30c",
   26299 => x"30c30c",
   26300 => x"30c30c",
   26301 => x"30c30c",
   26302 => x"30c32e",
   26303 => x"ffffff",
   26304 => x"ffffff",
   26305 => x"ffffff",
   26306 => x"ffffff",
   26307 => x"ffffff",
   26308 => x"ffffff",
   26309 => x"ffffff",
   26310 => x"fffa95",
   26311 => x"abffff",
   26312 => x"ffffff",
   26313 => x"ffffff",
   26314 => x"ffffff",
   26315 => x"ffffff",
   26316 => x"ffffff",
   26317 => x"ffffff",
   26318 => x"ffffff",
   26319 => x"ffffff",
   26320 => x"ffffff",
   26321 => x"fffeb0",
   26322 => x"c30c30",
   26323 => x"c30c30",
   26324 => x"c30c30",
   26325 => x"c30c30",
   26326 => x"c30c30",
   26327 => x"c30c30",
   26328 => x"c30c30",
   26329 => x"c30c30",
   26330 => x"c30c30",
   26331 => x"c30c30",
   26332 => x"c30c30",
   26333 => x"820820",
   26334 => x"820820",
   26335 => x"820820",
   26336 => x"820820",
   26337 => x"820820",
   26338 => x"820820",
   26339 => x"820820",
   26340 => x"820820",
   26341 => x"820820",
   26342 => x"820820",
   26343 => x"820820",
   26344 => x"820820",
   26345 => x"820820",
   26346 => x"820820",
   26347 => x"820820",
   26348 => x"820820",
   26349 => x"820820",
   26350 => x"820820",
   26351 => x"820820",
   26352 => x"820820",
   26353 => x"820820",
   26354 => x"820820",
   26355 => x"820410",
   26356 => x"410410",
   26357 => x"410410",
   26358 => x"410410",
   26359 => x"410410",
   26360 => x"410410",
   26361 => x"410410",
   26362 => x"410410",
   26363 => x"410410",
   26364 => x"410410",
   26365 => x"410410",
   26366 => x"410410",
   26367 => x"410410",
   26368 => x"410410",
   26369 => x"410410",
   26370 => x"410410",
   26371 => x"410410",
   26372 => x"410410",
   26373 => x"410410",
   26374 => x"410410",
   26375 => x"410410",
   26376 => x"410410",
   26377 => x"410410",
   26378 => x"410000",
   26379 => x"000000",
   26380 => x"000000",
   26381 => x"000000",
   26382 => x"000000",
   26383 => x"000000",
   26384 => x"000000",
   26385 => x"000000",
   26386 => x"000000",
   26387 => x"000000",
   26388 => x"000000",
   26389 => x"00057f",
   26390 => x"ffffff",
   26391 => x"ffffff",
   26392 => x"ffffff",
   26393 => x"ffffd5",
   26394 => x"00002a",
   26395 => x"ffffff",
   26396 => x"ffffff",
   26397 => x"fffa80",
   26398 => x"00002a",
   26399 => x"ffffff",
   26400 => x"ffffff",
   26401 => x"ffffff",
   26402 => x"ffffff",
   26403 => x"ffffff",
   26404 => x"ffffff",
   26405 => x"ffffff",
   26406 => x"d70c30",
   26407 => x"c30c30",
   26408 => x"c30c30",
   26409 => x"c30c30",
   26410 => x"c30c30",
   26411 => x"c30c30",
   26412 => x"867cf3",
   26413 => x"cf3cf3",
   26414 => x"cf3cf3",
   26415 => x"cf3cf3",
   26416 => x"cf3cf3",
   26417 => x"cf3cf3",
   26418 => x"cf3cf3",
   26419 => x"cf3cf3",
   26420 => x"cf3cf3",
   26421 => x"cf3cf3",
   26422 => x"cf3cf3",
   26423 => x"cf3cf3",
   26424 => x"cf3cf3",
   26425 => x"cf3cf3",
   26426 => x"cf3cf3",
   26427 => x"cf3dea",
   26428 => x"bbffff",
   26429 => x"ffffff",
   26430 => x"ffffff",
   26431 => x"ffffff",
   26432 => x"ffffff",
   26433 => x"ffffff",
   26434 => x"ffffff",
   26435 => x"ffffff",
   26436 => x"ffffff",
   26437 => x"ffffff",
   26438 => x"ffffff",
   26439 => x"ffffff",
   26440 => x"fee74e",
   26441 => x"3cf3cf",
   26442 => x"3cf3cf",
   26443 => x"3cf3cf",
   26444 => x"3cf3cf",
   26445 => x"3cf3cf",
   26446 => x"3cf3cf",
   26447 => x"3cf3cf",
   26448 => x"3cf3cf",
   26449 => x"3cf3cf",
   26450 => x"3cf3cf",
   26451 => x"3cf3cf",
   26452 => x"3cf3cf",
   26453 => x"3cf3cf",
   26454 => x"3cf3cf",
   26455 => x"3cf3cf",
   26456 => x"3cd30c",
   26457 => x"30c30c",
   26458 => x"30c30c",
   26459 => x"30c30c",
   26460 => x"30c30c",
   26461 => x"30c30c",
   26462 => x"30cbbf",
   26463 => x"ffffff",
   26464 => x"ffffff",
   26465 => x"ffffff",
   26466 => x"ffffff",
   26467 => x"ffffff",
   26468 => x"ffffff",
   26469 => x"ffffff",
   26470 => x"fea56a",
   26471 => x"ffffff",
   26472 => x"ffffff",
   26473 => x"ffffff",
   26474 => x"ffffff",
   26475 => x"ffffff",
   26476 => x"ffffff",
   26477 => x"ffffff",
   26478 => x"ffffff",
   26479 => x"ffffff",
   26480 => x"ffffff",
   26481 => x"fffeb0",
   26482 => x"c30c30",
   26483 => x"c30c30",
   26484 => x"c30c30",
   26485 => x"c30c30",
   26486 => x"c30c30",
   26487 => x"c30c30",
   26488 => x"c30c30",
   26489 => x"c30c30",
   26490 => x"c30c30",
   26491 => x"c30c30",
   26492 => x"c30c30",
   26493 => x"820820",
   26494 => x"820820",
   26495 => x"820820",
   26496 => x"820820",
   26497 => x"820820",
   26498 => x"820820",
   26499 => x"820820",
   26500 => x"820820",
   26501 => x"820820",
   26502 => x"820820",
   26503 => x"820820",
   26504 => x"820820",
   26505 => x"820820",
   26506 => x"820820",
   26507 => x"820820",
   26508 => x"820820",
   26509 => x"820820",
   26510 => x"820820",
   26511 => x"820820",
   26512 => x"820820",
   26513 => x"820820",
   26514 => x"820820",
   26515 => x"820410",
   26516 => x"410410",
   26517 => x"410410",
   26518 => x"410410",
   26519 => x"410410",
   26520 => x"410410",
   26521 => x"410410",
   26522 => x"410410",
   26523 => x"410410",
   26524 => x"410410",
   26525 => x"410410",
   26526 => x"410410",
   26527 => x"410410",
   26528 => x"410410",
   26529 => x"410410",
   26530 => x"410410",
   26531 => x"410410",
   26532 => x"410410",
   26533 => x"410410",
   26534 => x"410410",
   26535 => x"410410",
   26536 => x"410410",
   26537 => x"410410",
   26538 => x"410000",
   26539 => x"000000",
   26540 => x"000000",
   26541 => x"000000",
   26542 => x"000000",
   26543 => x"000000",
   26544 => x"000000",
   26545 => x"000000",
   26546 => x"000000",
   26547 => x"000000",
   26548 => x"000000",
   26549 => x"00057f",
   26550 => x"ffffff",
   26551 => x"ffffff",
   26552 => x"ffffff",
   26553 => x"ffffd5",
   26554 => x"00002a",
   26555 => x"ffffff",
   26556 => x"ffffff",
   26557 => x"ffffd5",
   26558 => x"000015",
   26559 => x"ffffff",
   26560 => x"ffffff",
   26561 => x"ffffff",
   26562 => x"ffffff",
   26563 => x"ffffff",
   26564 => x"ffffff",
   26565 => x"ffffff",
   26566 => x"ff5c30",
   26567 => x"c30c30",
   26568 => x"c30c30",
   26569 => x"c30c30",
   26570 => x"c30c30",
   26571 => x"c30c30",
   26572 => x"867cf3",
   26573 => x"cf3cf3",
   26574 => x"cf3cf3",
   26575 => x"cf3cf3",
   26576 => x"cf3cf3",
   26577 => x"cf3cf3",
   26578 => x"cf3cf3",
   26579 => x"cf3cf3",
   26580 => x"cf3cf3",
   26581 => x"cf3cf3",
   26582 => x"cf3cf3",
   26583 => x"cf3cf3",
   26584 => x"cf3cf3",
   26585 => x"cf3cf3",
   26586 => x"cf3cf3",
   26587 => x"cf3cf7",
   26588 => x"aaefff",
   26589 => x"ffffff",
   26590 => x"ffffff",
   26591 => x"ffffff",
   26592 => x"ffffff",
   26593 => x"ffffff",
   26594 => x"ffffff",
   26595 => x"ffffff",
   26596 => x"ffffff",
   26597 => x"ffffff",
   26598 => x"ffffff",
   26599 => x"ffffff",
   26600 => x"fdd38f",
   26601 => x"3cf3cf",
   26602 => x"3cf3cf",
   26603 => x"3cf3cf",
   26604 => x"3cf3cf",
   26605 => x"3cf3cf",
   26606 => x"3cf3cf",
   26607 => x"3cf3cf",
   26608 => x"3cf3cf",
   26609 => x"3cf3cf",
   26610 => x"3cf3cf",
   26611 => x"3cf3cf",
   26612 => x"3cf3cf",
   26613 => x"3cf3cf",
   26614 => x"3cf3cf",
   26615 => x"3cf3cf",
   26616 => x"3ce30c",
   26617 => x"30c30c",
   26618 => x"30c30c",
   26619 => x"30c30c",
   26620 => x"30c30c",
   26621 => x"30c30c",
   26622 => x"32efff",
   26623 => x"ffffff",
   26624 => x"ffffff",
   26625 => x"ffffff",
   26626 => x"ffffff",
   26627 => x"ffffff",
   26628 => x"ffffff",
   26629 => x"ffffff",
   26630 => x"a95abf",
   26631 => x"ffffff",
   26632 => x"ffffff",
   26633 => x"ffffff",
   26634 => x"ffffff",
   26635 => x"ffffff",
   26636 => x"ffffff",
   26637 => x"ffffff",
   26638 => x"ffffff",
   26639 => x"ffffff",
   26640 => x"ffffff",
   26641 => x"fffeb0",
   26642 => x"c30c30",
   26643 => x"c30c30",
   26644 => x"c30c30",
   26645 => x"c30c30",
   26646 => x"c30c30",
   26647 => x"c30c30",
   26648 => x"c30c30",
   26649 => x"c30c30",
   26650 => x"c30c30",
   26651 => x"c30c30",
   26652 => x"c30c30",
   26653 => x"820820",
   26654 => x"820820",
   26655 => x"820820",
   26656 => x"820820",
   26657 => x"820820",
   26658 => x"820820",
   26659 => x"820820",
   26660 => x"820820",
   26661 => x"820820",
   26662 => x"820820",
   26663 => x"820820",
   26664 => x"820820",
   26665 => x"820820",
   26666 => x"820820",
   26667 => x"820820",
   26668 => x"820820",
   26669 => x"820820",
   26670 => x"820820",
   26671 => x"820820",
   26672 => x"820820",
   26673 => x"820820",
   26674 => x"820820",
   26675 => x"820410",
   26676 => x"410410",
   26677 => x"410410",
   26678 => x"410410",
   26679 => x"410410",
   26680 => x"410410",
   26681 => x"410410",
   26682 => x"410410",
   26683 => x"410410",
   26684 => x"410410",
   26685 => x"410410",
   26686 => x"410410",
   26687 => x"410410",
   26688 => x"410410",
   26689 => x"410410",
   26690 => x"410410",
   26691 => x"410410",
   26692 => x"410410",
   26693 => x"410410",
   26694 => x"410410",
   26695 => x"410410",
   26696 => x"410410",
   26697 => x"410410",
   26698 => x"410000",
   26699 => x"000000",
   26700 => x"000000",
   26701 => x"000000",
   26702 => x"000000",
   26703 => x"000000",
   26704 => x"000000",
   26705 => x"000000",
   26706 => x"000000",
   26707 => x"000000",
   26708 => x"000000",
   26709 => x"00057f",
   26710 => x"ffffff",
   26711 => x"ffffff",
   26712 => x"ffffff",
   26713 => x"ffffd5",
   26714 => x"00002a",
   26715 => x"ffffff",
   26716 => x"ffffff",
   26717 => x"ffffea",
   26718 => x"000000",
   26719 => x"abffff",
   26720 => x"ffffff",
   26721 => x"ffffff",
   26722 => x"ffffff",
   26723 => x"ffffff",
   26724 => x"ffffff",
   26725 => x"ffffff",
   26726 => x"ffad70",
   26727 => x"c30c30",
   26728 => x"c30c30",
   26729 => x"c30c30",
   26730 => x"c30c30",
   26731 => x"c30c30",
   26732 => x"8b7cf3",
   26733 => x"cf3cf3",
   26734 => x"cf3cf3",
   26735 => x"cf3cf3",
   26736 => x"cf3cf3",
   26737 => x"cf3cf3",
   26738 => x"cf3cf3",
   26739 => x"cf3cf3",
   26740 => x"cf3cf3",
   26741 => x"cf3cf3",
   26742 => x"cf3cf3",
   26743 => x"cf3cf3",
   26744 => x"cf3cf3",
   26745 => x"cf3cf3",
   26746 => x"cf3cf3",
   26747 => x"cf3cf3",
   26748 => x"9eabbf",
   26749 => x"ffffff",
   26750 => x"ffffff",
   26751 => x"ffffff",
   26752 => x"ffffff",
   26753 => x"ffffff",
   26754 => x"ffffff",
   26755 => x"ffffff",
   26756 => x"ffffff",
   26757 => x"ffffff",
   26758 => x"ffffff",
   26759 => x"ffffff",
   26760 => x"74e3cf",
   26761 => x"3cf3cf",
   26762 => x"3cf3cf",
   26763 => x"3cf3cf",
   26764 => x"3cf3cf",
   26765 => x"3cf3cf",
   26766 => x"3cf3cf",
   26767 => x"3cf3cf",
   26768 => x"3cf3cf",
   26769 => x"3cf3cf",
   26770 => x"3cf3cf",
   26771 => x"3cf3cf",
   26772 => x"3cf3cf",
   26773 => x"3cf3cf",
   26774 => x"3cf3cf",
   26775 => x"3cf3cf",
   26776 => x"3ce30c",
   26777 => x"30c30c",
   26778 => x"30c30c",
   26779 => x"30c30c",
   26780 => x"30c30c",
   26781 => x"30c30c",
   26782 => x"bbffff",
   26783 => x"ffffff",
   26784 => x"ffffff",
   26785 => x"ffffff",
   26786 => x"ffffff",
   26787 => x"ffffff",
   26788 => x"ffffff",
   26789 => x"ffffea",
   26790 => x"56afff",
   26791 => x"ffffff",
   26792 => x"ffffff",
   26793 => x"ffffff",
   26794 => x"ffffff",
   26795 => x"ffffff",
   26796 => x"ffffff",
   26797 => x"ffffff",
   26798 => x"ffffff",
   26799 => x"ffffff",
   26800 => x"ffffff",
   26801 => x"fffeb0",
   26802 => x"c30c30",
   26803 => x"c30c30",
   26804 => x"c30c30",
   26805 => x"c30c30",
   26806 => x"c30c30",
   26807 => x"c30c30",
   26808 => x"c30c30",
   26809 => x"c30c30",
   26810 => x"c30c30",
   26811 => x"c30c30",
   26812 => x"c30c30",
   26813 => x"820820",
   26814 => x"820820",
   26815 => x"820820",
   26816 => x"820820",
   26817 => x"820820",
   26818 => x"820820",
   26819 => x"820820",
   26820 => x"820820",
   26821 => x"820820",
   26822 => x"820820",
   26823 => x"820820",
   26824 => x"820820",
   26825 => x"820820",
   26826 => x"820820",
   26827 => x"820820",
   26828 => x"820820",
   26829 => x"820820",
   26830 => x"820820",
   26831 => x"820820",
   26832 => x"820820",
   26833 => x"820820",
   26834 => x"820820",
   26835 => x"820410",
   26836 => x"410410",
   26837 => x"410410",
   26838 => x"410410",
   26839 => x"410410",
   26840 => x"410410",
   26841 => x"410410",
   26842 => x"410410",
   26843 => x"410410",
   26844 => x"410410",
   26845 => x"410410",
   26846 => x"410410",
   26847 => x"410410",
   26848 => x"410410",
   26849 => x"410410",
   26850 => x"410410",
   26851 => x"410410",
   26852 => x"410410",
   26853 => x"410410",
   26854 => x"410410",
   26855 => x"410410",
   26856 => x"410410",
   26857 => x"410410",
   26858 => x"410000",
   26859 => x"000000",
   26860 => x"000000",
   26861 => x"000000",
   26862 => x"000000",
   26863 => x"000000",
   26864 => x"000000",
   26865 => x"000000",
   26866 => x"000000",
   26867 => x"000000",
   26868 => x"000000",
   26869 => x"00057f",
   26870 => x"ffffff",
   26871 => x"ffffff",
   26872 => x"ffffff",
   26873 => x"ffffd5",
   26874 => x"00002a",
   26875 => x"ffffff",
   26876 => x"ffffff",
   26877 => x"ffffff",
   26878 => x"540000",
   26879 => x"57ffff",
   26880 => x"ffffff",
   26881 => x"ffffff",
   26882 => x"ffffff",
   26883 => x"ffffff",
   26884 => x"ffffff",
   26885 => x"ffffff",
   26886 => x"fffeb5",
   26887 => x"c30c30",
   26888 => x"c30c30",
   26889 => x"c30c30",
   26890 => x"c30c30",
   26891 => x"c30c31",
   26892 => x"5f7cf3",
   26893 => x"cf3cf3",
   26894 => x"cf3cf3",
   26895 => x"cf3cf3",
   26896 => x"cf3cf3",
   26897 => x"cf3cf3",
   26898 => x"cf3cf3",
   26899 => x"cf3cf3",
   26900 => x"cf3cf3",
   26901 => x"cf3cf3",
   26902 => x"cf3cf3",
   26903 => x"cf3cf3",
   26904 => x"cf3cf3",
   26905 => x"cf3cf3",
   26906 => x"cf3cf3",
   26907 => x"cf3cf3",
   26908 => x"ce7aae",
   26909 => x"ffffff",
   26910 => x"ffffff",
   26911 => x"ffffff",
   26912 => x"ffffff",
   26913 => x"ffffff",
   26914 => x"ffffff",
   26915 => x"ffffff",
   26916 => x"ffffff",
   26917 => x"ffffff",
   26918 => x"ffffff",
   26919 => x"ffffdd",
   26920 => x"34f3cf",
   26921 => x"3cf3cf",
   26922 => x"3cf3cf",
   26923 => x"3cf3cf",
   26924 => x"3cf3cf",
   26925 => x"3cf3cf",
   26926 => x"3cf3cf",
   26927 => x"3cf3cf",
   26928 => x"3cf3cf",
   26929 => x"3cf3cf",
   26930 => x"3cf3cf",
   26931 => x"3cf3cf",
   26932 => x"3cf3cf",
   26933 => x"3cf3cf",
   26934 => x"3cf3cf",
   26935 => x"3cf3cf",
   26936 => x"3ce34c",
   26937 => x"30c30c",
   26938 => x"30c30c",
   26939 => x"30c30c",
   26940 => x"30c30c",
   26941 => x"30c31d",
   26942 => x"ffffff",
   26943 => x"ffffff",
   26944 => x"ffffff",
   26945 => x"ffffff",
   26946 => x"ffffff",
   26947 => x"ffffff",
   26948 => x"ffffff",
   26949 => x"ffffd5",
   26950 => x"57ffff",
   26951 => x"ffffff",
   26952 => x"ffffff",
   26953 => x"ffffff",
   26954 => x"ffffff",
   26955 => x"ffffff",
   26956 => x"ffffff",
   26957 => x"ffffff",
   26958 => x"ffffff",
   26959 => x"ffffff",
   26960 => x"ffffff",
   26961 => x"fffeb0",
   26962 => x"c30c30",
   26963 => x"c30c30",
   26964 => x"c30c30",
   26965 => x"c30c30",
   26966 => x"c30c30",
   26967 => x"c30c30",
   26968 => x"c30c30",
   26969 => x"c30c30",
   26970 => x"c30c30",
   26971 => x"c30c30",
   26972 => x"c30c30",
   26973 => x"820820",
   26974 => x"820820",
   26975 => x"820820",
   26976 => x"820820",
   26977 => x"820820",
   26978 => x"820820",
   26979 => x"820820",
   26980 => x"820820",
   26981 => x"820820",
   26982 => x"820820",
   26983 => x"820820",
   26984 => x"820820",
   26985 => x"820820",
   26986 => x"820820",
   26987 => x"820820",
   26988 => x"820820",
   26989 => x"820820",
   26990 => x"820820",
   26991 => x"820820",
   26992 => x"820820",
   26993 => x"820820",
   26994 => x"820820",
   26995 => x"820410",
   26996 => x"410410",
   26997 => x"410410",
   26998 => x"410410",
   26999 => x"410410",
   27000 => x"410410",
   27001 => x"410410",
   27002 => x"410410",
   27003 => x"410410",
   27004 => x"410410",
   27005 => x"410410",
   27006 => x"410410",
   27007 => x"410410",
   27008 => x"410410",
   27009 => x"410410",
   27010 => x"410410",
   27011 => x"410410",
   27012 => x"410410",
   27013 => x"410410",
   27014 => x"410410",
   27015 => x"410410",
   27016 => x"410410",
   27017 => x"410410",
   27018 => x"410000",
   27019 => x"000000",
   27020 => x"000000",
   27021 => x"000000",
   27022 => x"000000",
   27023 => x"000000",
   27024 => x"000000",
   27025 => x"000000",
   27026 => x"000000",
   27027 => x"000000",
   27028 => x"000000",
   27029 => x"00057f",
   27030 => x"ffffff",
   27031 => x"ffffff",
   27032 => x"ffffff",
   27033 => x"ffffd5",
   27034 => x"00002a",
   27035 => x"ffffff",
   27036 => x"ffffff",
   27037 => x"ffffff",
   27038 => x"a80000",
   27039 => x"02afff",
   27040 => x"ffffff",
   27041 => x"ffffff",
   27042 => x"ffffff",
   27043 => x"ffffff",
   27044 => x"ffffff",
   27045 => x"ffffff",
   27046 => x"fffffa",
   27047 => x"d70c30",
   27048 => x"c30c30",
   27049 => x"c30c30",
   27050 => x"c30c30",
   27051 => x"c30c21",
   27052 => x"9f3cf3",
   27053 => x"cf3cf3",
   27054 => x"cf3cf3",
   27055 => x"cf3cf3",
   27056 => x"cf3cf3",
   27057 => x"cf3cf3",
   27058 => x"cf3cf3",
   27059 => x"cf3cf3",
   27060 => x"cf3cf3",
   27061 => x"cf3cf3",
   27062 => x"cf3cf3",
   27063 => x"cf3cf3",
   27064 => x"cf3cf3",
   27065 => x"cf3cf3",
   27066 => x"cf3cf3",
   27067 => x"cf3cf3",
   27068 => x"cf399a",
   27069 => x"bbffff",
   27070 => x"ffffff",
   27071 => x"ffffff",
   27072 => x"ffffff",
   27073 => x"ffffff",
   27074 => x"ffffff",
   27075 => x"ffffff",
   27076 => x"ffffff",
   27077 => x"ffffff",
   27078 => x"ffffff",
   27079 => x"fff74d",
   27080 => x"3cf3cf",
   27081 => x"3cf3cf",
   27082 => x"3cf3cf",
   27083 => x"3cf3cf",
   27084 => x"3cf3cf",
   27085 => x"3cf3cf",
   27086 => x"3cf3cf",
   27087 => x"3cf3cf",
   27088 => x"3cf3cf",
   27089 => x"3cf3cf",
   27090 => x"3cf3cf",
   27091 => x"3cf3cf",
   27092 => x"3cf3cf",
   27093 => x"3cf3cf",
   27094 => x"3cf3cf",
   27095 => x"3cf3cf",
   27096 => x"3cf34c",
   27097 => x"30c30c",
   27098 => x"30c30c",
   27099 => x"30c30c",
   27100 => x"30c30c",
   27101 => x"30c77f",
   27102 => x"ffffff",
   27103 => x"ffffff",
   27104 => x"ffffff",
   27105 => x"ffffff",
   27106 => x"ffffff",
   27107 => x"ffffff",
   27108 => x"ffffff",
   27109 => x"fffa95",
   27110 => x"abffff",
   27111 => x"ffffff",
   27112 => x"ffffff",
   27113 => x"ffffff",
   27114 => x"ffffff",
   27115 => x"ffffff",
   27116 => x"ffffff",
   27117 => x"ffffff",
   27118 => x"ffffff",
   27119 => x"ffffff",
   27120 => x"ffffff",
   27121 => x"fffeb0",
   27122 => x"c30c30",
   27123 => x"c30c30",
   27124 => x"c30c30",
   27125 => x"c30c30",
   27126 => x"c30c30",
   27127 => x"c30c30",
   27128 => x"c30c30",
   27129 => x"c30c30",
   27130 => x"c30c30",
   27131 => x"c30c30",
   27132 => x"c30c30",
   27133 => x"820820",
   27134 => x"820820",
   27135 => x"820820",
   27136 => x"820820",
   27137 => x"820820",
   27138 => x"820820",
   27139 => x"820820",
   27140 => x"820820",
   27141 => x"820820",
   27142 => x"820820",
   27143 => x"820820",
   27144 => x"820820",
   27145 => x"820820",
   27146 => x"820820",
   27147 => x"820820",
   27148 => x"820820",
   27149 => x"820820",
   27150 => x"820820",
   27151 => x"820820",
   27152 => x"820820",
   27153 => x"820820",
   27154 => x"820820",
   27155 => x"820410",
   27156 => x"410410",
   27157 => x"410410",
   27158 => x"410410",
   27159 => x"410410",
   27160 => x"410410",
   27161 => x"410410",
   27162 => x"410410",
   27163 => x"410410",
   27164 => x"410410",
   27165 => x"410410",
   27166 => x"410410",
   27167 => x"410410",
   27168 => x"410410",
   27169 => x"410410",
   27170 => x"410410",
   27171 => x"410410",
   27172 => x"410410",
   27173 => x"410410",
   27174 => x"410410",
   27175 => x"410410",
   27176 => x"410410",
   27177 => x"410410",
   27178 => x"410000",
   27179 => x"000000",
   27180 => x"000000",
   27181 => x"000000",
   27182 => x"000000",
   27183 => x"000000",
   27184 => x"000000",
   27185 => x"000000",
   27186 => x"000000",
   27187 => x"000000",
   27188 => x"000000",
   27189 => x"00057f",
   27190 => x"ffffff",
   27191 => x"ffffff",
   27192 => x"ffffff",
   27193 => x"ffffd5",
   27194 => x"00002a",
   27195 => x"ffffff",
   27196 => x"ffffff",
   27197 => x"ffffff",
   27198 => x"fd5000",
   27199 => x"015fff",
   27200 => x"ffffff",
   27201 => x"ffffff",
   27202 => x"ffffff",
   27203 => x"ffffff",
   27204 => x"ffffff",
   27205 => x"ffffff",
   27206 => x"ffffff",
   27207 => x"eb5c30",
   27208 => x"c30c30",
   27209 => x"c30c30",
   27210 => x"c30c30",
   27211 => x"c30c21",
   27212 => x"9f3cf3",
   27213 => x"cf3cf3",
   27214 => x"cf3cf3",
   27215 => x"cf3cf3",
   27216 => x"cf3cf3",
   27217 => x"cf3cf3",
   27218 => x"cf3cf3",
   27219 => x"cf3cf3",
   27220 => x"cf3cf3",
   27221 => x"cf3cf3",
   27222 => x"cf3cf3",
   27223 => x"cf3cf3",
   27224 => x"cf3cf3",
   27225 => x"cf3cf3",
   27226 => x"cf3cf3",
   27227 => x"cf3cf3",
   27228 => x"cf3ce6",
   27229 => x"6aefff",
   27230 => x"ffffff",
   27231 => x"ffffff",
   27232 => x"ffffff",
   27233 => x"ffffff",
   27234 => x"ffffff",
   27235 => x"ffffff",
   27236 => x"ffffff",
   27237 => x"ffffff",
   27238 => x"ffffff",
   27239 => x"fdd34f",
   27240 => x"3cf3cf",
   27241 => x"3cf3cf",
   27242 => x"3cf3cf",
   27243 => x"3cf3cf",
   27244 => x"3cf3cf",
   27245 => x"3cf3cf",
   27246 => x"3cf3cf",
   27247 => x"3cf3cf",
   27248 => x"3cf3cf",
   27249 => x"3cf3cf",
   27250 => x"3cf3cf",
   27251 => x"3cf3cf",
   27252 => x"3cf3cf",
   27253 => x"3cf3cf",
   27254 => x"3cf3cf",
   27255 => x"3cf3cf",
   27256 => x"3cf38c",
   27257 => x"30c30c",
   27258 => x"30c30c",
   27259 => x"30c30c",
   27260 => x"30c30c",
   27261 => x"31dfff",
   27262 => x"ffffff",
   27263 => x"ffffff",
   27264 => x"ffffff",
   27265 => x"ffffff",
   27266 => x"ffffff",
   27267 => x"ffffff",
   27268 => x"ffffff",
   27269 => x"fffa95",
   27270 => x"abffff",
   27271 => x"ffffff",
   27272 => x"ffffff",
   27273 => x"ffffff",
   27274 => x"ffffff",
   27275 => x"ffffff",
   27276 => x"ffffff",
   27277 => x"ffffff",
   27278 => x"ffffff",
   27279 => x"ffffff",
   27280 => x"ffffff",
   27281 => x"fffeb0",
   27282 => x"c30c30",
   27283 => x"c30c30",
   27284 => x"c30c30",
   27285 => x"c30c30",
   27286 => x"c30c30",
   27287 => x"c30c30",
   27288 => x"c30c30",
   27289 => x"c30c30",
   27290 => x"c30c30",
   27291 => x"c30c30",
   27292 => x"c30c30",
   27293 => x"820820",
   27294 => x"820820",
   27295 => x"820820",
   27296 => x"820820",
   27297 => x"820820",
   27298 => x"820820",
   27299 => x"820820",
   27300 => x"820820",
   27301 => x"820820",
   27302 => x"820820",
   27303 => x"820820",
   27304 => x"820820",
   27305 => x"820820",
   27306 => x"820820",
   27307 => x"820820",
   27308 => x"820820",
   27309 => x"820820",
   27310 => x"820820",
   27311 => x"820820",
   27312 => x"820820",
   27313 => x"820820",
   27314 => x"820820",
   27315 => x"820410",
   27316 => x"410410",
   27317 => x"410410",
   27318 => x"410410",
   27319 => x"410410",
   27320 => x"410410",
   27321 => x"410410",
   27322 => x"410410",
   27323 => x"410410",
   27324 => x"410410",
   27325 => x"410410",
   27326 => x"410410",
   27327 => x"410410",
   27328 => x"410410",
   27329 => x"410410",
   27330 => x"410410",
   27331 => x"410410",
   27332 => x"410410",
   27333 => x"410410",
   27334 => x"410410",
   27335 => x"410410",
   27336 => x"410410",
   27337 => x"410410",
   27338 => x"410000",
   27339 => x"000000",
   27340 => x"000000",
   27341 => x"000000",
   27342 => x"000000",
   27343 => x"000000",
   27344 => x"000000",
   27345 => x"000000",
   27346 => x"000000",
   27347 => x"000000",
   27348 => x"000000",
   27349 => x"00057f",
   27350 => x"ffffff",
   27351 => x"ffffff",
   27352 => x"ffffff",
   27353 => x"ffffd5",
   27354 => x"00002a",
   27355 => x"ffffff",
   27356 => x"ffffff",
   27357 => x"ffffff",
   27358 => x"fea000",
   27359 => x"000abf",
   27360 => x"ffffff",
   27361 => x"ffffff",
   27362 => x"ffffff",
   27363 => x"ffffff",
   27364 => x"ffffff",
   27365 => x"ffffff",
   27366 => x"ffffff",
   27367 => x"ffad70",
   27368 => x"c30c30",
   27369 => x"c30c30",
   27370 => x"c30c30",
   27371 => x"c30c22",
   27372 => x"df3cf3",
   27373 => x"cf3cf3",
   27374 => x"cf3cf3",
   27375 => x"cf3cf3",
   27376 => x"cf3cf3",
   27377 => x"cf3cf3",
   27378 => x"cf3cf3",
   27379 => x"cf3cf3",
   27380 => x"cf3cf3",
   27381 => x"cf3cf3",
   27382 => x"cf3cf3",
   27383 => x"cf3cf3",
   27384 => x"cf3cf3",
   27385 => x"cf3cf3",
   27386 => x"cf3cf3",
   27387 => x"cf3cf3",
   27388 => x"cf3cf3",
   27389 => x"99abbf",
   27390 => x"ffffff",
   27391 => x"ffffff",
   27392 => x"ffffff",
   27393 => x"ffffff",
   27394 => x"ffffff",
   27395 => x"ffffff",
   27396 => x"ffffff",
   27397 => x"ffffff",
   27398 => x"ffffee",
   27399 => x"74e3cf",
   27400 => x"3cf3cf",
   27401 => x"3cf3cf",
   27402 => x"3cf3cf",
   27403 => x"3cf3cf",
   27404 => x"3cf3cf",
   27405 => x"3cf3cf",
   27406 => x"3cf3cf",
   27407 => x"3cf3cf",
   27408 => x"3cf3cf",
   27409 => x"3cf3cf",
   27410 => x"3cf3cf",
   27411 => x"3cf3cf",
   27412 => x"3cf3cf",
   27413 => x"3cf3cf",
   27414 => x"3cf3cf",
   27415 => x"3cf3cf",
   27416 => x"3cf38c",
   27417 => x"30c30c",
   27418 => x"30c30c",
   27419 => x"30c30c",
   27420 => x"30c30c",
   27421 => x"77ffff",
   27422 => x"ffffff",
   27423 => x"ffffff",
   27424 => x"ffffff",
   27425 => x"ffffff",
   27426 => x"ffffff",
   27427 => x"ffffff",
   27428 => x"ffffff",
   27429 => x"fffa95",
   27430 => x"abffff",
   27431 => x"ffffff",
   27432 => x"ffffff",
   27433 => x"ffffff",
   27434 => x"ffffff",
   27435 => x"ffffff",
   27436 => x"ffffff",
   27437 => x"ffffff",
   27438 => x"ffffff",
   27439 => x"ffffff",
   27440 => x"ffffff",
   27441 => x"fffeb0",
   27442 => x"c30c30",
   27443 => x"c30c30",
   27444 => x"c30c30",
   27445 => x"c30c30",
   27446 => x"c30c30",
   27447 => x"c30c30",
   27448 => x"c30c30",
   27449 => x"c30c30",
   27450 => x"c30c30",
   27451 => x"c30c30",
   27452 => x"c30c30",
   27453 => x"820820",
   27454 => x"820820",
   27455 => x"820820",
   27456 => x"820820",
   27457 => x"820820",
   27458 => x"820820",
   27459 => x"820820",
   27460 => x"820820",
   27461 => x"820820",
   27462 => x"820820",
   27463 => x"820820",
   27464 => x"820820",
   27465 => x"820820",
   27466 => x"820820",
   27467 => x"820820",
   27468 => x"820820",
   27469 => x"820820",
   27470 => x"820820",
   27471 => x"820820",
   27472 => x"820820",
   27473 => x"820820",
   27474 => x"820820",
   27475 => x"820410",
   27476 => x"410410",
   27477 => x"410410",
   27478 => x"410410",
   27479 => x"410410",
   27480 => x"410410",
   27481 => x"410410",
   27482 => x"410410",
   27483 => x"410410",
   27484 => x"410410",
   27485 => x"410410",
   27486 => x"410410",
   27487 => x"410410",
   27488 => x"410410",
   27489 => x"410410",
   27490 => x"410410",
   27491 => x"410410",
   27492 => x"410410",
   27493 => x"410410",
   27494 => x"410410",
   27495 => x"410410",
   27496 => x"410410",
   27497 => x"410410",
   27498 => x"410000",
   27499 => x"000000",
   27500 => x"000000",
   27501 => x"000000",
   27502 => x"000000",
   27503 => x"000000",
   27504 => x"000000",
   27505 => x"000000",
   27506 => x"000000",
   27507 => x"000000",
   27508 => x"000000",
   27509 => x"00057f",
   27510 => x"ffffff",
   27511 => x"ffffff",
   27512 => x"ffffff",
   27513 => x"ffffd5",
   27514 => x"55556a",
   27515 => x"ffffff",
   27516 => x"ffffff",
   27517 => x"ffffff",
   27518 => x"fff555",
   27519 => x"555abf",
   27520 => x"ffffff",
   27521 => x"ffffff",
   27522 => x"ffffff",
   27523 => x"ffffff",
   27524 => x"ffffff",
   27525 => x"ffffff",
   27526 => x"ffffff",
   27527 => x"fffeb5",
   27528 => x"c30c30",
   27529 => x"c30c30",
   27530 => x"c30c30",
   27531 => x"c30857",
   27532 => x"df3cf3",
   27533 => x"cf3cf3",
   27534 => x"cf3cf3",
   27535 => x"cf3cf3",
   27536 => x"cf3cf3",
   27537 => x"cf3cf3",
   27538 => x"cf3cf3",
   27539 => x"cf3cf3",
   27540 => x"cf3cf3",
   27541 => x"cf3cf3",
   27542 => x"cf3cf3",
   27543 => x"cf3cf3",
   27544 => x"cf3cf3",
   27545 => x"cf3cf3",
   27546 => x"cf3cf3",
   27547 => x"cf3cf3",
   27548 => x"cf3cf3",
   27549 => x"ce7aae",
   27550 => x"ffffff",
   27551 => x"ffffff",
   27552 => x"ffffff",
   27553 => x"ffffff",
   27554 => x"ffffff",
   27555 => x"ffffff",
   27556 => x"ffffff",
   27557 => x"ffffff",
   27558 => x"fffb9d",
   27559 => x"38f3cf",
   27560 => x"3cf3cf",
   27561 => x"3cf3cf",
   27562 => x"3cf3cf",
   27563 => x"3cf3cf",
   27564 => x"3cf3cf",
   27565 => x"3cf3cf",
   27566 => x"3cf3cf",
   27567 => x"3cf3cf",
   27568 => x"3cf3cf",
   27569 => x"3cf3cf",
   27570 => x"3cf3cf",
   27571 => x"3cf3cf",
   27572 => x"3cf3cf",
   27573 => x"3cf3cf",
   27574 => x"3cf3cf",
   27575 => x"3cf3cf",
   27576 => x"3cf38d",
   27577 => x"30c30c",
   27578 => x"30c30c",
   27579 => x"30c30c",
   27580 => x"30c31d",
   27581 => x"ffffff",
   27582 => x"ffffff",
   27583 => x"ffffff",
   27584 => x"ffffff",
   27585 => x"ffffff",
   27586 => x"ffffff",
   27587 => x"ffffff",
   27588 => x"ffffff",
   27589 => x"fffa95",
   27590 => x"abffff",
   27591 => x"ffffff",
   27592 => x"ffffff",
   27593 => x"ffffff",
   27594 => x"ffffff",
   27595 => x"ffffff",
   27596 => x"ffffff",
   27597 => x"ffffff",
   27598 => x"ffffff",
   27599 => x"ffffff",
   27600 => x"ffffff",
   27601 => x"fffeb0",
   27602 => x"c30c30",
   27603 => x"c30c30",
   27604 => x"c30c30",
   27605 => x"c30c30",
   27606 => x"c30c30",
   27607 => x"c30c30",
   27608 => x"c30c30",
   27609 => x"c30c30",
   27610 => x"c30c30",
   27611 => x"c30c30",
   27612 => x"c30c30",
   27613 => x"820820",
   27614 => x"820820",
   27615 => x"820820",
   27616 => x"820820",
   27617 => x"820820",
   27618 => x"820820",
   27619 => x"820820",
   27620 => x"820820",
   27621 => x"820820",
   27622 => x"820820",
   27623 => x"820820",
   27624 => x"820820",
   27625 => x"820820",
   27626 => x"820820",
   27627 => x"820820",
   27628 => x"820820",
   27629 => x"820820",
   27630 => x"820820",
   27631 => x"820820",
   27632 => x"820820",
   27633 => x"820820",
   27634 => x"820820",
   27635 => x"820410",
   27636 => x"410410",
   27637 => x"410410",
   27638 => x"410410",
   27639 => x"410410",
   27640 => x"410410",
   27641 => x"410410",
   27642 => x"410410",
   27643 => x"410410",
   27644 => x"410410",
   27645 => x"410410",
   27646 => x"410410",
   27647 => x"410410",
   27648 => x"410410",
   27649 => x"410410",
   27650 => x"410410",
   27651 => x"410410",
   27652 => x"410410",
   27653 => x"410410",
   27654 => x"410410",
   27655 => x"410410",
   27656 => x"410410",
   27657 => x"410410",
   27658 => x"410000",
   27659 => x"000000",
   27660 => x"000000",
   27661 => x"000000",
   27662 => x"000000",
   27663 => x"000000",
   27664 => x"000000",
   27665 => x"000000",
   27666 => x"000000",
   27667 => x"000000",
   27668 => x"000000",
   27669 => x"00057f",
   27670 => x"ffffff",
   27671 => x"ffffff",
   27672 => x"ffffff",
   27673 => x"ffffea",
   27674 => x"aaaabf",
   27675 => x"ffffff",
   27676 => x"ffffff",
   27677 => x"ffffff",
   27678 => x"ffffea",
   27679 => x"aaaabf",
   27680 => x"ffffff",
   27681 => x"ffffff",
   27682 => x"ffffff",
   27683 => x"ffffff",
   27684 => x"ffffff",
   27685 => x"ffffff",
   27686 => x"ffffff",
   27687 => x"fffffa",
   27688 => x"d70c30",
   27689 => x"c30c30",
   27690 => x"c30c30",
   27691 => x"c30867",
   27692 => x"cf3cf3",
   27693 => x"cf3cf3",
   27694 => x"cf3cf3",
   27695 => x"cf3cf3",
   27696 => x"cf3cf3",
   27697 => x"cf3cf3",
   27698 => x"cf3cf3",
   27699 => x"cf3cf3",
   27700 => x"cf3cf3",
   27701 => x"cf3cf3",
   27702 => x"cf3cf3",
   27703 => x"cf3cf3",
   27704 => x"cf3cf3",
   27705 => x"cf3cf3",
   27706 => x"cf3cf3",
   27707 => x"cf3cf3",
   27708 => x"cf3cf3",
   27709 => x"cf39ea",
   27710 => x"bbffff",
   27711 => x"ffffff",
   27712 => x"ffffff",
   27713 => x"ffffff",
   27714 => x"ffffff",
   27715 => x"ffffff",
   27716 => x"ffffff",
   27717 => x"ffffff",
   27718 => x"fee74e",
   27719 => x"3cf3cf",
   27720 => x"3cf3cf",
   27721 => x"3cf3cf",
   27722 => x"3cf3cf",
   27723 => x"3cf3cf",
   27724 => x"3cf3cf",
   27725 => x"3cf3cf",
   27726 => x"3cf3cf",
   27727 => x"3cf3cf",
   27728 => x"3cf3cf",
   27729 => x"3cf3cf",
   27730 => x"3cf3cf",
   27731 => x"3cf3cf",
   27732 => x"3cf3cf",
   27733 => x"3cf3cf",
   27734 => x"3cf3cf",
   27735 => x"3cf3cf",
   27736 => x"3cf3cd",
   27737 => x"30c30c",
   27738 => x"30c30c",
   27739 => x"30c30c",
   27740 => x"30cbbf",
   27741 => x"ffffff",
   27742 => x"ffffff",
   27743 => x"ffffff",
   27744 => x"ffffff",
   27745 => x"ffffff",
   27746 => x"ffffff",
   27747 => x"ffffff",
   27748 => x"ffffff",
   27749 => x"fffa95",
   27750 => x"abffff",
   27751 => x"ffffff",
   27752 => x"ffffff",
   27753 => x"ffffff",
   27754 => x"ffffff",
   27755 => x"ffffff",
   27756 => x"ffffff",
   27757 => x"ffffff",
   27758 => x"ffffff",
   27759 => x"ffffff",
   27760 => x"ffffff",
   27761 => x"fffeb0",
   27762 => x"c30c30",
   27763 => x"c30c30",
   27764 => x"c30c30",
   27765 => x"c30c30",
   27766 => x"c30c30",
   27767 => x"c30c30",
   27768 => x"c30c30",
   27769 => x"c30c30",
   27770 => x"c30c30",
   27771 => x"c30c30",
   27772 => x"c30c30",
   27773 => x"820820",
   27774 => x"820820",
   27775 => x"820820",
   27776 => x"820820",
   27777 => x"820820",
   27778 => x"820820",
   27779 => x"820820",
   27780 => x"820820",
   27781 => x"820820",
   27782 => x"820820",
   27783 => x"820820",
   27784 => x"820820",
   27785 => x"820820",
   27786 => x"820820",
   27787 => x"820820",
   27788 => x"820820",
   27789 => x"820820",
   27790 => x"820820",
   27791 => x"820820",
   27792 => x"820820",
   27793 => x"820820",
   27794 => x"820820",
   27795 => x"820410",
   27796 => x"410410",
   27797 => x"410410",
   27798 => x"410410",
   27799 => x"410410",
   27800 => x"410410",
   27801 => x"410410",
   27802 => x"410410",
   27803 => x"410410",
   27804 => x"410410",
   27805 => x"410410",
   27806 => x"410410",
   27807 => x"410410",
   27808 => x"410410",
   27809 => x"410410",
   27810 => x"410410",
   27811 => x"410410",
   27812 => x"410410",
   27813 => x"410410",
   27814 => x"410410",
   27815 => x"410410",
   27816 => x"410410",
   27817 => x"410410",
   27818 => x"410000",
   27819 => x"000000",
   27820 => x"000000",
   27821 => x"000000",
   27822 => x"000000",
   27823 => x"000000",
   27824 => x"000000",
   27825 => x"000000",
   27826 => x"000000",
   27827 => x"000000",
   27828 => x"000000",
   27829 => x"00057f",
   27830 => x"ffffff",
   27831 => x"ffffff",
   27832 => x"ffffff",
   27833 => x"ffffff",
   27834 => x"ffffff",
   27835 => x"ffffff",
   27836 => x"ffffff",
   27837 => x"ffffff",
   27838 => x"ffffff",
   27839 => x"ffffff",
   27840 => x"ffffff",
   27841 => x"ffffff",
   27842 => x"ffffff",
   27843 => x"ffffff",
   27844 => x"ffffff",
   27845 => x"ffffff",
   27846 => x"ffffff",
   27847 => x"ffffff",
   27848 => x"ff5c30",
   27849 => x"c30c30",
   27850 => x"c30c30",
   27851 => x"c30867",
   27852 => x"cf3cf3",
   27853 => x"cf3cf3",
   27854 => x"cf3cf3",
   27855 => x"cf3cf3",
   27856 => x"cf3cf3",
   27857 => x"cf3cf3",
   27858 => x"cf3cf3",
   27859 => x"cf3cf3",
   27860 => x"cf3cf3",
   27861 => x"cf3cf3",
   27862 => x"cf3cf3",
   27863 => x"cf3cf3",
   27864 => x"cf3cf3",
   27865 => x"cf3cf3",
   27866 => x"cf3cf3",
   27867 => x"cf3cf3",
   27868 => x"cf3cf3",
   27869 => x"cf3ce7",
   27870 => x"aaefff",
   27871 => x"ffffff",
   27872 => x"ffffff",
   27873 => x"ffffff",
   27874 => x"ffffff",
   27875 => x"ffffff",
   27876 => x"ffffff",
   27877 => x"ffffff",
   27878 => x"b9d38f",
   27879 => x"3cf3cf",
   27880 => x"3cf3cf",
   27881 => x"3cf3cf",
   27882 => x"3cf3cf",
   27883 => x"3cf3cf",
   27884 => x"3cf3cf",
   27885 => x"3cf3cf",
   27886 => x"3cf3cf",
   27887 => x"3cf3cf",
   27888 => x"3cf3cf",
   27889 => x"3cf3cf",
   27890 => x"3cf3cf",
   27891 => x"3cf3cf",
   27892 => x"3cf3cf",
   27893 => x"3cf3cf",
   27894 => x"3cf3cf",
   27895 => x"3cf3cf",
   27896 => x"3cf3ce",
   27897 => x"30c30c",
   27898 => x"30c30c",
   27899 => x"30c30c",
   27900 => x"32efff",
   27901 => x"ffffff",
   27902 => x"ffffff",
   27903 => x"ffffff",
   27904 => x"ffffff",
   27905 => x"ffffff",
   27906 => x"ffffff",
   27907 => x"ffffff",
   27908 => x"ffffff",
   27909 => x"fffa95",
   27910 => x"abffff",
   27911 => x"ffffff",
   27912 => x"ffffff",
   27913 => x"ffffff",
   27914 => x"ffffff",
   27915 => x"ffffff",
   27916 => x"ffffff",
   27917 => x"ffffff",
   27918 => x"ffffff",
   27919 => x"ffffff",
   27920 => x"ffffff",
   27921 => x"fffeb0",
   27922 => x"c30c30",
   27923 => x"c30c30",
   27924 => x"c30c30",
   27925 => x"c30c30",
   27926 => x"c30c30",
   27927 => x"c30c30",
   27928 => x"c30c30",
   27929 => x"c30c30",
   27930 => x"c30c30",
   27931 => x"c30c30",
   27932 => x"c30c30",
   27933 => x"820820",
   27934 => x"820820",
   27935 => x"820820",
   27936 => x"820820",
   27937 => x"820820",
   27938 => x"820820",
   27939 => x"820820",
   27940 => x"820820",
   27941 => x"820820",
   27942 => x"820820",
   27943 => x"820820",
   27944 => x"820820",
   27945 => x"820820",
   27946 => x"820820",
   27947 => x"820820",
   27948 => x"820820",
   27949 => x"820820",
   27950 => x"820820",
   27951 => x"820820",
   27952 => x"820820",
   27953 => x"820820",
   27954 => x"820820",
   27955 => x"820410",
   27956 => x"410410",
   27957 => x"410410",
   27958 => x"410410",
   27959 => x"410410",
   27960 => x"410410",
   27961 => x"410410",
   27962 => x"410410",
   27963 => x"410410",
   27964 => x"410410",
   27965 => x"410410",
   27966 => x"410410",
   27967 => x"410410",
   27968 => x"410410",
   27969 => x"410410",
   27970 => x"410410",
   27971 => x"410410",
   27972 => x"410410",
   27973 => x"410410",
   27974 => x"410410",
   27975 => x"410410",
   27976 => x"410410",
   27977 => x"410410",
   27978 => x"410000",
   27979 => x"000000",
   27980 => x"000000",
   27981 => x"000000",
   27982 => x"000000",
   27983 => x"000000",
   27984 => x"000000",
   27985 => x"000000",
   27986 => x"000000",
   27987 => x"000000",
   27988 => x"000000",
   27989 => x"00057f",
   27990 => x"ffffff",
   27991 => x"ffffff",
   27992 => x"ffffff",
   27993 => x"ffffff",
   27994 => x"ffffff",
   27995 => x"ffffff",
   27996 => x"ffffff",
   27997 => x"ffffff",
   27998 => x"ffffff",
   27999 => x"ffffff",
   28000 => x"ffffff",
   28001 => x"ffffff",
   28002 => x"ffffff",
   28003 => x"ffffff",
   28004 => x"ffffff",
   28005 => x"ffffff",
   28006 => x"ffffff",
   28007 => x"ffffff",
   28008 => x"fffd70",
   28009 => x"c30c30",
   28010 => x"c30c30",
   28011 => x"c308b7",
   28012 => x"cf3cf3",
   28013 => x"cf3cf3",
   28014 => x"cf3cf3",
   28015 => x"cf3cf3",
   28016 => x"cf3cf3",
   28017 => x"cf3cf3",
   28018 => x"cf3cf3",
   28019 => x"cf3cf3",
   28020 => x"cf3cf3",
   28021 => x"cf3cf3",
   28022 => x"cf3cf3",
   28023 => x"cf3cf3",
   28024 => x"cf3cf3",
   28025 => x"cf3cf3",
   28026 => x"cf3cf3",
   28027 => x"cf3cf3",
   28028 => x"cf3cf3",
   28029 => x"cf3cf3",
   28030 => x"deabbf",
   28031 => x"ffffff",
   28032 => x"ffffff",
   28033 => x"ffffff",
   28034 => x"ffffff",
   28035 => x"ffffff",
   28036 => x"ffffff",
   28037 => x"ffffee",
   28038 => x"74e3cf",
   28039 => x"3cf3cf",
   28040 => x"3cf3cf",
   28041 => x"3cf3cf",
   28042 => x"3cf3cf",
   28043 => x"3cf3cf",
   28044 => x"3cf3cf",
   28045 => x"3cf3cf",
   28046 => x"3cf3cf",
   28047 => x"3cf3cf",
   28048 => x"3cf3cf",
   28049 => x"3cf3cf",
   28050 => x"3cf3cf",
   28051 => x"3cf3cf",
   28052 => x"3cf3cf",
   28053 => x"3cf3cf",
   28054 => x"3cf3cf",
   28055 => x"3cf3cf",
   28056 => x"3cf3ce",
   28057 => x"30c30c",
   28058 => x"30c30c",
   28059 => x"30c31d",
   28060 => x"bbffff",
   28061 => x"ffffff",
   28062 => x"ffffff",
   28063 => x"ffffff",
   28064 => x"ffffff",
   28065 => x"ffffff",
   28066 => x"ffffff",
   28067 => x"ffffff",
   28068 => x"ffffff",
   28069 => x"fffa95",
   28070 => x"abffff",
   28071 => x"ffffff",
   28072 => x"ffffff",
   28073 => x"ffffff",
   28074 => x"ffffff",
   28075 => x"ffffff",
   28076 => x"ffffff",
   28077 => x"ffffff",
   28078 => x"ffffff",
   28079 => x"ffffff",
   28080 => x"ffffff",
   28081 => x"fffeb0",
   28082 => x"c30c30",
   28083 => x"c30c30",
   28084 => x"c30c30",
   28085 => x"c30c30",
   28086 => x"c30c30",
   28087 => x"c30c30",
   28088 => x"c30c30",
   28089 => x"c30c30",
   28090 => x"c30c30",
   28091 => x"c30c30",
   28092 => x"c30c30",
   28093 => x"820820",
   28094 => x"820820",
   28095 => x"820820",
   28096 => x"820820",
   28097 => x"820820",
   28098 => x"820820",
   28099 => x"820820",
   28100 => x"820820",
   28101 => x"820820",
   28102 => x"820820",
   28103 => x"820820",
   28104 => x"820820",
   28105 => x"820820",
   28106 => x"820820",
   28107 => x"820820",
   28108 => x"820820",
   28109 => x"820820",
   28110 => x"820820",
   28111 => x"820820",
   28112 => x"820820",
   28113 => x"820820",
   28114 => x"820820",
   28115 => x"820410",
   28116 => x"410410",
   28117 => x"410410",
   28118 => x"410410",
   28119 => x"410410",
   28120 => x"410410",
   28121 => x"410410",
   28122 => x"410410",
   28123 => x"410410",
   28124 => x"410410",
   28125 => x"410410",
   28126 => x"410410",
   28127 => x"410410",
   28128 => x"410410",
   28129 => x"410410",
   28130 => x"410410",
   28131 => x"410410",
   28132 => x"410410",
   28133 => x"410410",
   28134 => x"410410",
   28135 => x"410410",
   28136 => x"410410",
   28137 => x"410410",
   28138 => x"410000",
   28139 => x"000000",
   28140 => x"000000",
   28141 => x"000000",
   28142 => x"000000",
   28143 => x"000000",
   28144 => x"000000",
   28145 => x"000000",
   28146 => x"000000",
   28147 => x"000000",
   28148 => x"000000",
   28149 => x"00057f",
   28150 => x"ffffff",
   28151 => x"ffffff",
   28152 => x"ffffff",
   28153 => x"ffffff",
   28154 => x"ffffff",
   28155 => x"ffffff",
   28156 => x"ffffff",
   28157 => x"ffffff",
   28158 => x"ffffff",
   28159 => x"ffffff",
   28160 => x"ffffff",
   28161 => x"ffffff",
   28162 => x"ffffff",
   28163 => x"ffffff",
   28164 => x"ffffff",
   28165 => x"ffffff",
   28166 => x"ffffff",
   28167 => x"ffffff",
   28168 => x"fffffa",
   28169 => x"d70c30",
   28170 => x"c30c30",
   28171 => x"c309b7",
   28172 => x"cf3cf3",
   28173 => x"cf3cf3",
   28174 => x"cf3cf3",
   28175 => x"cf3cf3",
   28176 => x"cf3cf3",
   28177 => x"cf3cf3",
   28178 => x"cf3cf3",
   28179 => x"cf3cf3",
   28180 => x"cf3cf3",
   28181 => x"cf3cf3",
   28182 => x"cf3cf3",
   28183 => x"cf3cf3",
   28184 => x"cf3cf3",
   28185 => x"cf3cf3",
   28186 => x"cf3cf3",
   28187 => x"cf3cf3",
   28188 => x"cf3cf3",
   28189 => x"cf3cf3",
   28190 => x"cf399e",
   28191 => x"bfffff",
   28192 => x"ffffff",
   28193 => x"ffffff",
   28194 => x"ffffff",
   28195 => x"ffffff",
   28196 => x"ffffff",
   28197 => x"fffb9d",
   28198 => x"38f3cf",
   28199 => x"3cf3cf",
   28200 => x"3cf3cf",
   28201 => x"3cf3cf",
   28202 => x"3cf3cf",
   28203 => x"3cf3cf",
   28204 => x"3cf3cf",
   28205 => x"3cf3cf",
   28206 => x"3cf3cf",
   28207 => x"3cf3cf",
   28208 => x"3cf3cf",
   28209 => x"3cf3cf",
   28210 => x"3cf3cf",
   28211 => x"3cf3cf",
   28212 => x"3cf3cf",
   28213 => x"3cf3cf",
   28214 => x"3cf3cf",
   28215 => x"3cf3cf",
   28216 => x"3cf3ce",
   28217 => x"30c30c",
   28218 => x"30c30c",
   28219 => x"30c76e",
   28220 => x"ffffff",
   28221 => x"ffffff",
   28222 => x"ffffff",
   28223 => x"ffffff",
   28224 => x"ffffff",
   28225 => x"ffffff",
   28226 => x"ffffff",
   28227 => x"ffffff",
   28228 => x"ffffff",
   28229 => x"fffa95",
   28230 => x"abffff",
   28231 => x"ffffff",
   28232 => x"ffffff",
   28233 => x"ffffff",
   28234 => x"ffffff",
   28235 => x"ffffff",
   28236 => x"ffffff",
   28237 => x"ffffff",
   28238 => x"ffffff",
   28239 => x"ffffff",
   28240 => x"ffffff",
   28241 => x"fffeb0",
   28242 => x"c30c30",
   28243 => x"c30c30",
   28244 => x"c30c30",
   28245 => x"c30c30",
   28246 => x"c30c30",
   28247 => x"c30c30",
   28248 => x"c30c30",
   28249 => x"c30c30",
   28250 => x"c30c30",
   28251 => x"c30c30",
   28252 => x"c30c30",
   28253 => x"820820",
   28254 => x"820820",
   28255 => x"820820",
   28256 => x"820820",
   28257 => x"820820",
   28258 => x"820820",
   28259 => x"820820",
   28260 => x"820820",
   28261 => x"820820",
   28262 => x"820820",
   28263 => x"820820",
   28264 => x"820820",
   28265 => x"820820",
   28266 => x"820820",
   28267 => x"820820",
   28268 => x"820820",
   28269 => x"820820",
   28270 => x"820820",
   28271 => x"820820",
   28272 => x"820820",
   28273 => x"820820",
   28274 => x"820820",
   28275 => x"820410",
   28276 => x"410410",
   28277 => x"410410",
   28278 => x"410410",
   28279 => x"410410",
   28280 => x"410410",
   28281 => x"410410",
   28282 => x"410410",
   28283 => x"410410",
   28284 => x"410410",
   28285 => x"410410",
   28286 => x"410410",
   28287 => x"410410",
   28288 => x"410410",
   28289 => x"410410",
   28290 => x"410410",
   28291 => x"410410",
   28292 => x"410410",
   28293 => x"410410",
   28294 => x"410410",
   28295 => x"410410",
   28296 => x"410410",
   28297 => x"410410",
   28298 => x"410000",
   28299 => x"000000",
   28300 => x"000000",
   28301 => x"000000",
   28302 => x"000000",
   28303 => x"000000",
   28304 => x"000000",
   28305 => x"000000",
   28306 => x"000000",
   28307 => x"000000",
   28308 => x"000000",
   28309 => x"00057f",
   28310 => x"ffffff",
   28311 => x"ffffff",
   28312 => x"ffffff",
   28313 => x"ffffff",
   28314 => x"ffffff",
   28315 => x"ffffff",
   28316 => x"ffffff",
   28317 => x"ffffff",
   28318 => x"ffffff",
   28319 => x"ffffff",
   28320 => x"ffffff",
   28321 => x"ffffff",
   28322 => x"ffffff",
   28323 => x"ffffff",
   28324 => x"ffffff",
   28325 => x"ffffff",
   28326 => x"ffffff",
   28327 => x"ffffff",
   28328 => x"ffffff",
   28329 => x"eb5c30",
   28330 => x"c30c30",
   28331 => x"c319b7",
   28332 => x"cf3cf3",
   28333 => x"cf3cf3",
   28334 => x"cf3cf3",
   28335 => x"cf3cf3",
   28336 => x"cf3cf3",
   28337 => x"cf3cf3",
   28338 => x"cf3cf3",
   28339 => x"cf3cf3",
   28340 => x"cf3cf3",
   28341 => x"cf3cf3",
   28342 => x"cf3cf3",
   28343 => x"cf3cf3",
   28344 => x"cf3cf3",
   28345 => x"cf3cf3",
   28346 => x"cf3cf3",
   28347 => x"cf3cf3",
   28348 => x"cf3cf3",
   28349 => x"cf3cf3",
   28350 => x"cf3ce6",
   28351 => x"6aefff",
   28352 => x"ffffff",
   28353 => x"ffffff",
   28354 => x"ffffff",
   28355 => x"ffffff",
   28356 => x"ffffff",
   28357 => x"fde34e",
   28358 => x"3cf3cf",
   28359 => x"3cf3cf",
   28360 => x"3cf3cf",
   28361 => x"3cf3cf",
   28362 => x"3cf3cf",
   28363 => x"3cf3cf",
   28364 => x"3cf3cf",
   28365 => x"3cf3cf",
   28366 => x"3cf3cf",
   28367 => x"3cf3cf",
   28368 => x"3cf3cf",
   28369 => x"3cf3cf",
   28370 => x"3cf3cf",
   28371 => x"3cf3cf",
   28372 => x"3cf3cf",
   28373 => x"3cf3cf",
   28374 => x"3cf3cf",
   28375 => x"3cf3cf",
   28376 => x"3cf3ce",
   28377 => x"34c30c",
   28378 => x"30c30c",
   28379 => x"31dfff",
   28380 => x"ffffff",
   28381 => x"ffffff",
   28382 => x"ffffff",
   28383 => x"ffffff",
   28384 => x"ffffff",
   28385 => x"ffffff",
   28386 => x"ffffff",
   28387 => x"ffffff",
   28388 => x"ffffff",
   28389 => x"fffa95",
   28390 => x"abffff",
   28391 => x"ffffff",
   28392 => x"ffffff",
   28393 => x"ffffff",
   28394 => x"ffffff",
   28395 => x"ffffff",
   28396 => x"ffffff",
   28397 => x"ffffff",
   28398 => x"ffffff",
   28399 => x"ffffff",
   28400 => x"ffffff",
   28401 => x"fffeb0",
   28402 => x"c30c30",
   28403 => x"c30c30",
   28404 => x"c30c30",
   28405 => x"c30c30",
   28406 => x"c30c30",
   28407 => x"c30c30",
   28408 => x"c30c30",
   28409 => x"c30c30",
   28410 => x"c30c30",
   28411 => x"c30c30",
   28412 => x"c30c30",
   28413 => x"820820",
   28414 => x"820820",
   28415 => x"820820",
   28416 => x"820820",
   28417 => x"820820",
   28418 => x"820820",
   28419 => x"820820",
   28420 => x"820820",
   28421 => x"820820",
   28422 => x"820820",
   28423 => x"820820",
   28424 => x"820820",
   28425 => x"820820",
   28426 => x"820820",
   28427 => x"820820",
   28428 => x"820820",
   28429 => x"820820",
   28430 => x"820820",
   28431 => x"820820",
   28432 => x"820820",
   28433 => x"820820",
   28434 => x"820820",
   28435 => x"820410",
   28436 => x"410410",
   28437 => x"410410",
   28438 => x"410410",
   28439 => x"410410",
   28440 => x"410410",
   28441 => x"410410",
   28442 => x"410410",
   28443 => x"410410",
   28444 => x"410410",
   28445 => x"410410",
   28446 => x"410410",
   28447 => x"410410",
   28448 => x"410410",
   28449 => x"410410",
   28450 => x"410410",
   28451 => x"410410",
   28452 => x"410410",
   28453 => x"410410",
   28454 => x"410410",
   28455 => x"410410",
   28456 => x"410410",
   28457 => x"410410",
   28458 => x"410000",
   28459 => x"000000",
   28460 => x"000000",
   28461 => x"000000",
   28462 => x"000000",
   28463 => x"000000",
   28464 => x"000000",
   28465 => x"000000",
   28466 => x"000000",
   28467 => x"000000",
   28468 => x"000000",
   28469 => x"00057f",
   28470 => x"ffffff",
   28471 => x"ffffff",
   28472 => x"ffffff",
   28473 => x"ffffff",
   28474 => x"ffffff",
   28475 => x"ffffff",
   28476 => x"ffffff",
   28477 => x"ffffff",
   28478 => x"ffffff",
   28479 => x"ffffff",
   28480 => x"ffffff",
   28481 => x"ffffff",
   28482 => x"ffffff",
   28483 => x"ffffff",
   28484 => x"ffffff",
   28485 => x"ffffff",
   28486 => x"ffffff",
   28487 => x"ffffff",
   28488 => x"ffffff",
   28489 => x"ffad70",
   28490 => x"c30c30",
   28491 => x"c319f3",
   28492 => x"cf3cf3",
   28493 => x"cf3cf3",
   28494 => x"cf3cf3",
   28495 => x"cf3cf3",
   28496 => x"cf3cf3",
   28497 => x"cf3cf3",
   28498 => x"cf3cf3",
   28499 => x"cf3cf3",
   28500 => x"cf3cf3",
   28501 => x"cf3cf3",
   28502 => x"cf3cf3",
   28503 => x"cf3cf3",
   28504 => x"cf3cf3",
   28505 => x"cf3cf3",
   28506 => x"cf3cf3",
   28507 => x"cf3cf3",
   28508 => x"cf3cf3",
   28509 => x"cf3cf3",
   28510 => x"cf3cf3",
   28511 => x"9dabbf",
   28512 => x"ffffff",
   28513 => x"ffffff",
   28514 => x"ffffff",
   28515 => x"ffffff",
   28516 => x"ffffee",
   28517 => x"78e3cf",
   28518 => x"3cf3cf",
   28519 => x"3cf3cf",
   28520 => x"3cf3cf",
   28521 => x"3cf3cf",
   28522 => x"3cf3cf",
   28523 => x"3cf3cf",
   28524 => x"3cf3cf",
   28525 => x"3cf3cf",
   28526 => x"3cf3cf",
   28527 => x"3cf3cf",
   28528 => x"3cf3cf",
   28529 => x"3cf3cf",
   28530 => x"3cf3cf",
   28531 => x"3cf3cf",
   28532 => x"3cf3cf",
   28533 => x"3cf3cf",
   28534 => x"3cf3cf",
   28535 => x"3cf3cf",
   28536 => x"3cf3cf",
   28537 => x"34c30c",
   28538 => x"30c31d",
   28539 => x"bbffff",
   28540 => x"ffffff",
   28541 => x"ffffff",
   28542 => x"ffffff",
   28543 => x"ffffff",
   28544 => x"ffffff",
   28545 => x"ffffff",
   28546 => x"ffffff",
   28547 => x"ffffff",
   28548 => x"ffffff",
   28549 => x"fffa95",
   28550 => x"abffff",
   28551 => x"ffffff",
   28552 => x"ffffff",
   28553 => x"ffffff",
   28554 => x"ffffff",
   28555 => x"ffffff",
   28556 => x"ffffff",
   28557 => x"ffffff",
   28558 => x"ffffff",
   28559 => x"ffffff",
   28560 => x"ffffff",
   28561 => x"fffeb0",
   28562 => x"c30c30",
   28563 => x"c30c30",
   28564 => x"c30c30",
   28565 => x"c30c30",
   28566 => x"c30c30",
   28567 => x"c30c30",
   28568 => x"c30c30",
   28569 => x"c30c30",
   28570 => x"c30c30",
   28571 => x"c30c30",
   28572 => x"c30c30",
   28573 => x"820820",
   28574 => x"820820",
   28575 => x"820820",
   28576 => x"820820",
   28577 => x"820820",
   28578 => x"820820",
   28579 => x"820820",
   28580 => x"820820",
   28581 => x"820820",
   28582 => x"820820",
   28583 => x"820820",
   28584 => x"820820",
   28585 => x"820820",
   28586 => x"820820",
   28587 => x"820820",
   28588 => x"820820",
   28589 => x"820820",
   28590 => x"820820",
   28591 => x"820820",
   28592 => x"820820",
   28593 => x"820820",
   28594 => x"820820",
   28595 => x"820410",
   28596 => x"410410",
   28597 => x"410410",
   28598 => x"410410",
   28599 => x"410410",
   28600 => x"410410",
   28601 => x"410410",
   28602 => x"410410",
   28603 => x"410410",
   28604 => x"410410",
   28605 => x"410410",
   28606 => x"410410",
   28607 => x"410410",
   28608 => x"410410",
   28609 => x"410410",
   28610 => x"410410",
   28611 => x"410410",
   28612 => x"410410",
   28613 => x"410410",
   28614 => x"410410",
   28615 => x"410410",
   28616 => x"410410",
   28617 => x"410410",
   28618 => x"410000",
   28619 => x"000000",
   28620 => x"000000",
   28621 => x"000000",
   28622 => x"000000",
   28623 => x"000000",
   28624 => x"000000",
   28625 => x"000000",
   28626 => x"000000",
   28627 => x"000000",
   28628 => x"000000",
   28629 => x"00057f",
   28630 => x"ffffff",
   28631 => x"ffffff",
   28632 => x"ffffff",
   28633 => x"ffffff",
   28634 => x"ffffff",
   28635 => x"ffffff",
   28636 => x"ffffff",
   28637 => x"ffffff",
   28638 => x"ffffff",
   28639 => x"ffffff",
   28640 => x"ffffff",
   28641 => x"ffffff",
   28642 => x"ffffff",
   28643 => x"ffffff",
   28644 => x"ffffff",
   28645 => x"ffffff",
   28646 => x"ffffff",
   28647 => x"ffffff",
   28648 => x"ffffff",
   28649 => x"fffffa",
   28650 => x"c30c30",
   28651 => x"c319f3",
   28652 => x"cf3cf3",
   28653 => x"cf3cf3",
   28654 => x"cf3cf3",
   28655 => x"cf3cf3",
   28656 => x"cf3cf3",
   28657 => x"cf3cf3",
   28658 => x"cf3cf3",
   28659 => x"cf3cf3",
   28660 => x"cf3cf3",
   28661 => x"cf3cf3",
   28662 => x"cf3cf3",
   28663 => x"cf3cf3",
   28664 => x"cf3cf3",
   28665 => x"cf3cf3",
   28666 => x"cf3cf3",
   28667 => x"cf3cf3",
   28668 => x"cf3cf3",
   28669 => x"cf3cf3",
   28670 => x"cf3cf3",
   28671 => x"cf39ae",
   28672 => x"ffffff",
   28673 => x"ffffff",
   28674 => x"ffffff",
   28675 => x"ffffff",
   28676 => x"fffb9e",
   28677 => x"38f3cf",
   28678 => x"3cf3cf",
   28679 => x"3cf3cf",
   28680 => x"3cf3cf",
   28681 => x"3cf3cf",
   28682 => x"3cf3cf",
   28683 => x"3cf3cf",
   28684 => x"3cf3cf",
   28685 => x"3cf3cf",
   28686 => x"3cf3cf",
   28687 => x"3cf3cf",
   28688 => x"3cf3cf",
   28689 => x"3cf3cf",
   28690 => x"3cf3cf",
   28691 => x"3cf3cf",
   28692 => x"3cf3cf",
   28693 => x"3cf3cf",
   28694 => x"3cf3cf",
   28695 => x"3cf3cf",
   28696 => x"3cf3cf",
   28697 => x"34c30c",
   28698 => x"30c76e",
   28699 => x"ffffff",
   28700 => x"ffffff",
   28701 => x"ffffff",
   28702 => x"ffffff",
   28703 => x"ffffff",
   28704 => x"ffffff",
   28705 => x"ffffff",
   28706 => x"ffffff",
   28707 => x"ffffff",
   28708 => x"ffffff",
   28709 => x"fffa95",
   28710 => x"abffff",
   28711 => x"ffffff",
   28712 => x"ffffff",
   28713 => x"ffffff",
   28714 => x"ffffff",
   28715 => x"ffffff",
   28716 => x"ffffff",
   28717 => x"ffffff",
   28718 => x"ffffff",
   28719 => x"ffffff",
   28720 => x"ffffff",
   28721 => x"fffeb0",
   28722 => x"c30c30",
   28723 => x"c30c30",
   28724 => x"c30c30",
   28725 => x"c30c30",
   28726 => x"c30c30",
   28727 => x"c30c30",
   28728 => x"c30c30",
   28729 => x"c30c30",
   28730 => x"c30c30",
   28731 => x"c30c30",
   28732 => x"c30c30",
   28733 => x"820820",
   28734 => x"820820",
   28735 => x"820820",
   28736 => x"820820",
   28737 => x"820820",
   28738 => x"820820",
   28739 => x"820820",
   28740 => x"820820",
   28741 => x"820820",
   28742 => x"820820",
   28743 => x"820820",
   28744 => x"820820",
   28745 => x"820820",
   28746 => x"820820",
   28747 => x"820820",
   28748 => x"820820",
   28749 => x"820820",
   28750 => x"820820",
   28751 => x"820820",
   28752 => x"820820",
   28753 => x"820820",
   28754 => x"820820",
   28755 => x"820410",
   28756 => x"410410",
   28757 => x"410410",
   28758 => x"410410",
   28759 => x"410410",
   28760 => x"410410",
   28761 => x"410410",
   28762 => x"410410",
   28763 => x"410410",
   28764 => x"410410",
   28765 => x"410410",
   28766 => x"410410",
   28767 => x"410410",
   28768 => x"410410",
   28769 => x"410410",
   28770 => x"410410",
   28771 => x"410410",
   28772 => x"410410",
   28773 => x"410410",
   28774 => x"410410",
   28775 => x"410410",
   28776 => x"410410",
   28777 => x"410410",
   28778 => x"410000",
   28779 => x"000000",
   28780 => x"000000",
   28781 => x"000000",
   28782 => x"000000",
   28783 => x"000000",
   28784 => x"000000",
   28785 => x"000000",
   28786 => x"000000",
   28787 => x"000000",
   28788 => x"000000",
   28789 => x"00057f",
   28790 => x"ffffff",
   28791 => x"ffffff",
   28792 => x"ffffff",
   28793 => x"ffffff",
   28794 => x"ffffff",
   28795 => x"ffffff",
   28796 => x"ffffff",
   28797 => x"ffffff",
   28798 => x"ffffff",
   28799 => x"ffffff",
   28800 => x"ffffff",
   28801 => x"ffffff",
   28802 => x"ffffff",
   28803 => x"ffffff",
   28804 => x"ffffff",
   28805 => x"ffffff",
   28806 => x"ffffff",
   28807 => x"ffffff",
   28808 => x"ffffff",
   28809 => x"ffffff",
   28810 => x"eb5c30",
   28811 => x"c219f3",
   28812 => x"cf3cf3",
   28813 => x"cf3cf3",
   28814 => x"cf3cf3",
   28815 => x"cf3cf3",
   28816 => x"cf3cf3",
   28817 => x"cf3cf3",
   28818 => x"cf3cf3",
   28819 => x"cf3cf3",
   28820 => x"cf3cf3",
   28821 => x"cf3cf3",
   28822 => x"cf3cf3",
   28823 => x"cf3cf3",
   28824 => x"cf3cf3",
   28825 => x"cf3cf3",
   28826 => x"cf3cf3",
   28827 => x"cf3cf3",
   28828 => x"cf3cf3",
   28829 => x"cf3cf3",
   28830 => x"cf3cf3",
   28831 => x"cf3ce7",
   28832 => x"6aefff",
   28833 => x"ffffff",
   28834 => x"ffffff",
   28835 => x"ffffff",
   28836 => x"fee38f",
   28837 => x"3cf3cf",
   28838 => x"3cf3cf",
   28839 => x"3cf3cf",
   28840 => x"3cf3cf",
   28841 => x"3cf3cf",
   28842 => x"3cf3cf",
   28843 => x"3cf3cf",
   28844 => x"3cf3cf",
   28845 => x"3cf3cf",
   28846 => x"3cf3cf",
   28847 => x"3cf3cf",
   28848 => x"3cf3cf",
   28849 => x"3cf3cf",
   28850 => x"3cf3cf",
   28851 => x"3cf3cf",
   28852 => x"3cf3cf",
   28853 => x"3cf3cf",
   28854 => x"3cf3cf",
   28855 => x"3cf3cf",
   28856 => x"3cf3cf",
   28857 => x"38c30c",
   28858 => x"31dfff",
   28859 => x"ffffff",
   28860 => x"ffffff",
   28861 => x"ffffff",
   28862 => x"ffffff",
   28863 => x"ffffff",
   28864 => x"ffffff",
   28865 => x"ffffff",
   28866 => x"ffffff",
   28867 => x"ffffff",
   28868 => x"ffffff",
   28869 => x"fffa95",
   28870 => x"abffff",
   28871 => x"ffffff",
   28872 => x"ffffff",
   28873 => x"ffffff",
   28874 => x"ffffff",
   28875 => x"ffffff",
   28876 => x"ffffff",
   28877 => x"ffffff",
   28878 => x"ffffff",
   28879 => x"ffffff",
   28880 => x"ffffff",
   28881 => x"fffeb0",
   28882 => x"c30c30",
   28883 => x"c30c30",
   28884 => x"c30c30",
   28885 => x"c30c30",
   28886 => x"c30c30",
   28887 => x"c30c30",
   28888 => x"c30c30",
   28889 => x"c30c30",
   28890 => x"c30c30",
   28891 => x"c30c30",
   28892 => x"c30c30",
   28893 => x"820820",
   28894 => x"820820",
   28895 => x"820820",
   28896 => x"820820",
   28897 => x"820820",
   28898 => x"820820",
   28899 => x"820820",
   28900 => x"820820",
   28901 => x"820820",
   28902 => x"820820",
   28903 => x"820820",
   28904 => x"820820",
   28905 => x"820820",
   28906 => x"820820",
   28907 => x"820820",
   28908 => x"820820",
   28909 => x"820820",
   28910 => x"820820",
   28911 => x"820820",
   28912 => x"820820",
   28913 => x"820820",
   28914 => x"820820",
   28915 => x"820410",
   28916 => x"410410",
   28917 => x"410410",
   28918 => x"410410",
   28919 => x"410410",
   28920 => x"410410",
   28921 => x"410410",
   28922 => x"410410",
   28923 => x"410410",
   28924 => x"410410",
   28925 => x"410410",
   28926 => x"410410",
   28927 => x"410410",
   28928 => x"410410",
   28929 => x"410410",
   28930 => x"410410",
   28931 => x"410410",
   28932 => x"410410",
   28933 => x"410410",
   28934 => x"410410",
   28935 => x"410410",
   28936 => x"410410",
   28937 => x"410410",
   28938 => x"410000",
   28939 => x"000000",
   28940 => x"000000",
   28941 => x"000000",
   28942 => x"000000",
   28943 => x"000000",
   28944 => x"000000",
   28945 => x"000000",
   28946 => x"000000",
   28947 => x"000000",
   28948 => x"000000",
   28949 => x"00057f",
   28950 => x"ffffff",
   28951 => x"ffffff",
   28952 => x"ffffff",
   28953 => x"ffffff",
   28954 => x"ffffff",
   28955 => x"ffffff",
   28956 => x"ffffff",
   28957 => x"ffffff",
   28958 => x"ffffff",
   28959 => x"ffffff",
   28960 => x"ffffff",
   28961 => x"ffffff",
   28962 => x"ffffff",
   28963 => x"ffffff",
   28964 => x"ffffff",
   28965 => x"ffffff",
   28966 => x"ffffff",
   28967 => x"ffffff",
   28968 => x"ffffff",
   28969 => x"ffffff",
   28970 => x"fffd70",
   28971 => x"c219f3",
   28972 => x"cf3cf3",
   28973 => x"cf3cf3",
   28974 => x"cf3cf3",
   28975 => x"cf3cf3",
   28976 => x"cf3cf3",
   28977 => x"cf3cf3",
   28978 => x"cf3cf3",
   28979 => x"cf3cf3",
   28980 => x"cf3cf3",
   28981 => x"cf3cf3",
   28982 => x"cf3cf3",
   28983 => x"cf3cf3",
   28984 => x"cf3cf3",
   28985 => x"cf3cf3",
   28986 => x"cf3cf3",
   28987 => x"cf3cf3",
   28988 => x"cf3cf3",
   28989 => x"cf3cf3",
   28990 => x"cf3cf3",
   28991 => x"cf3cf3",
   28992 => x"ddabbf",
   28993 => x"ffffff",
   28994 => x"ffffff",
   28995 => x"ffffef",
   28996 => x"78e3cf",
   28997 => x"3cf3cf",
   28998 => x"3cf3cf",
   28999 => x"3cf3cf",
   29000 => x"3cf3cf",
   29001 => x"3cf3cf",
   29002 => x"3cf3cf",
   29003 => x"3cf3cf",
   29004 => x"3cf3cf",
   29005 => x"3cf3cf",
   29006 => x"3cf3cf",
   29007 => x"3cf3cf",
   29008 => x"3cf3cf",
   29009 => x"3cf3cf",
   29010 => x"3cf3cf",
   29011 => x"3cf3cf",
   29012 => x"3cf3cf",
   29013 => x"3cf3cf",
   29014 => x"3cf3cf",
   29015 => x"3cf3cf",
   29016 => x"3cf3cf",
   29017 => x"38c31d",
   29018 => x"bbffff",
   29019 => x"ffffff",
   29020 => x"ffffff",
   29021 => x"ffffff",
   29022 => x"ffffff",
   29023 => x"ffffff",
   29024 => x"ffffff",
   29025 => x"ffffff",
   29026 => x"ffffff",
   29027 => x"ffffff",
   29028 => x"ffffff",
   29029 => x"fffa95",
   29030 => x"abffff",
   29031 => x"ffffff",
   29032 => x"ffffff",
   29033 => x"ffffff",
   29034 => x"ffffff",
   29035 => x"ffffff",
   29036 => x"ffffff",
   29037 => x"ffffff",
   29038 => x"ffffff",
   29039 => x"ffffff",
   29040 => x"ffffff",
   29041 => x"fffeb0",
   29042 => x"c30c30",
   29043 => x"c30c30",
   29044 => x"c30c30",
   29045 => x"c30c30",
   29046 => x"c30c30",
   29047 => x"c30c30",
   29048 => x"c30c30",
   29049 => x"c30c30",
   29050 => x"c30c30",
   29051 => x"c30c30",
   29052 => x"c30c30",
   29053 => x"820820",
   29054 => x"820820",
   29055 => x"820820",
   29056 => x"820820",
   29057 => x"820820",
   29058 => x"820820",
   29059 => x"820820",
   29060 => x"820820",
   29061 => x"820820",
   29062 => x"820820",
   29063 => x"820820",
   29064 => x"820820",
   29065 => x"820820",
   29066 => x"820820",
   29067 => x"820820",
   29068 => x"820820",
   29069 => x"820820",
   29070 => x"820820",
   29071 => x"820820",
   29072 => x"820820",
   29073 => x"820820",
   29074 => x"820820",
   29075 => x"820410",
   29076 => x"410410",
   29077 => x"410410",
   29078 => x"410410",
   29079 => x"410410",
   29080 => x"410410",
   29081 => x"410410",
   29082 => x"410410",
   29083 => x"410410",
   29084 => x"410410",
   29085 => x"410410",
   29086 => x"410410",
   29087 => x"410410",
   29088 => x"410410",
   29089 => x"410410",
   29090 => x"410410",
   29091 => x"410410",
   29092 => x"410410",
   29093 => x"410410",
   29094 => x"410410",
   29095 => x"410410",
   29096 => x"410410",
   29097 => x"410410",
   29098 => x"410000",
   29099 => x"000000",
   29100 => x"000000",
   29101 => x"000000",
   29102 => x"000000",
   29103 => x"000000",
   29104 => x"000000",
   29105 => x"000000",
   29106 => x"000000",
   29107 => x"000000",
   29108 => x"000000",
   29109 => x"00057f",
   29110 => x"ffffff",
   29111 => x"ffffff",
   29112 => x"ffffff",
   29113 => x"ffffff",
   29114 => x"ffffff",
   29115 => x"ffffff",
   29116 => x"ffffff",
   29117 => x"ffffff",
   29118 => x"ffffff",
   29119 => x"ffffff",
   29120 => x"ffffff",
   29121 => x"ffffff",
   29122 => x"ffffff",
   29123 => x"ffffff",
   29124 => x"ffffff",
   29125 => x"ffffff",
   29126 => x"ffffff",
   29127 => x"ffffff",
   29128 => x"ffffff",
   29129 => x"ffffff",
   29130 => x"fffffa",
   29131 => x"d629f3",
   29132 => x"cf3cf3",
   29133 => x"cf3cf3",
   29134 => x"cf3cf3",
   29135 => x"cf3cf3",
   29136 => x"cf3cf3",
   29137 => x"cf3cf3",
   29138 => x"cf3cf3",
   29139 => x"cf3cf3",
   29140 => x"cf3cf3",
   29141 => x"cf3cf3",
   29142 => x"cf3cf3",
   29143 => x"cf3cf3",
   29144 => x"cf3cf3",
   29145 => x"cf3cf3",
   29146 => x"cf3cf3",
   29147 => x"cf3cf3",
   29148 => x"cf3cf3",
   29149 => x"cf3cf3",
   29150 => x"cf3cf3",
   29151 => x"cf3cf3",
   29152 => x"cf79da",
   29153 => x"bbffff",
   29154 => x"ffffff",
   29155 => x"fffb9e",
   29156 => x"3cf3cf",
   29157 => x"3cf3cf",
   29158 => x"3cf3cf",
   29159 => x"3cf3cf",
   29160 => x"3cf3cf",
   29161 => x"3cf3cf",
   29162 => x"3cf3cf",
   29163 => x"3cf3cf",
   29164 => x"3cf3cf",
   29165 => x"3cf3cf",
   29166 => x"3cf3cf",
   29167 => x"3cf3cf",
   29168 => x"3cf3cf",
   29169 => x"3cf3cf",
   29170 => x"3cf3cf",
   29171 => x"3cf3cf",
   29172 => x"3cf3cf",
   29173 => x"3cf3cf",
   29174 => x"3cf3cf",
   29175 => x"3cf3cf",
   29176 => x"3cf3cf",
   29177 => x"34c77f",
   29178 => x"ffffff",
   29179 => x"ffffff",
   29180 => x"ffffff",
   29181 => x"ffffff",
   29182 => x"ffffff",
   29183 => x"ffffff",
   29184 => x"ffffff",
   29185 => x"ffffff",
   29186 => x"ffffff",
   29187 => x"ffffff",
   29188 => x"ffffff",
   29189 => x"fffa95",
   29190 => x"abffff",
   29191 => x"ffffff",
   29192 => x"ffffff",
   29193 => x"ffffff",
   29194 => x"ffffff",
   29195 => x"ffffff",
   29196 => x"ffffff",
   29197 => x"ffffff",
   29198 => x"ffffff",
   29199 => x"ffffff",
   29200 => x"ffffff",
   29201 => x"fffeb0",
   29202 => x"c30c30",
   29203 => x"c30c30",
   29204 => x"c30c30",
   29205 => x"c30c30",
   29206 => x"c30c30",
   29207 => x"c30c30",
   29208 => x"c30c30",
   29209 => x"c30c30",
   29210 => x"c30c30",
   29211 => x"c30c30",
   29212 => x"c30c30",
   29213 => x"820820",
   29214 => x"820820",
   29215 => x"820820",
   29216 => x"820820",
   29217 => x"820820",
   29218 => x"820820",
   29219 => x"820820",
   29220 => x"820820",
   29221 => x"820820",
   29222 => x"820820",
   29223 => x"820820",
   29224 => x"820820",
   29225 => x"820820",
   29226 => x"820820",
   29227 => x"820820",
   29228 => x"820820",
   29229 => x"820820",
   29230 => x"820820",
   29231 => x"820820",
   29232 => x"820820",
   29233 => x"820820",
   29234 => x"820820",
   29235 => x"820410",
   29236 => x"410410",
   29237 => x"410410",
   29238 => x"410410",
   29239 => x"410410",
   29240 => x"410410",
   29241 => x"410410",
   29242 => x"410410",
   29243 => x"410410",
   29244 => x"410410",
   29245 => x"410410",
   29246 => x"410410",
   29247 => x"410410",
   29248 => x"410410",
   29249 => x"410410",
   29250 => x"410410",
   29251 => x"410410",
   29252 => x"410410",
   29253 => x"410410",
   29254 => x"410410",
   29255 => x"410410",
   29256 => x"410410",
   29257 => x"410410",
   29258 => x"410000",
   29259 => x"000000",
   29260 => x"000000",
   29261 => x"000000",
   29262 => x"000000",
   29263 => x"000000",
   29264 => x"000000",
   29265 => x"000000",
   29266 => x"000000",
   29267 => x"000000",
   29268 => x"000000",
   29269 => x"00057f",
   29270 => x"ffffff",
   29271 => x"ffffff",
   29272 => x"ffffff",
   29273 => x"ffffff",
   29274 => x"ffffff",
   29275 => x"ffffff",
   29276 => x"ffffff",
   29277 => x"ffffff",
   29278 => x"ffffff",
   29279 => x"ffffff",
   29280 => x"ffffff",
   29281 => x"ffffff",
   29282 => x"ffffff",
   29283 => x"ffffff",
   29284 => x"ffffff",
   29285 => x"ffffff",
   29286 => x"ffffff",
   29287 => x"ffffff",
   29288 => x"ffffff",
   29289 => x"ffffff",
   29290 => x"ffffff",
   29291 => x"ed75fb",
   29292 => x"df3cf3",
   29293 => x"cf3cf3",
   29294 => x"cf3cf3",
   29295 => x"cf3cf3",
   29296 => x"cf3cf3",
   29297 => x"cf3cf3",
   29298 => x"cf3cf3",
   29299 => x"cf3cf3",
   29300 => x"cf3cf3",
   29301 => x"cf3cf3",
   29302 => x"cf3cf3",
   29303 => x"cf3cf3",
   29304 => x"cf3cf3",
   29305 => x"cf3cf3",
   29306 => x"cf3cf3",
   29307 => x"cf3cf3",
   29308 => x"cf3cf3",
   29309 => x"cf3cf3",
   29310 => x"cf3cf3",
   29311 => x"cf3cf3",
   29312 => x"cf3cf7",
   29313 => x"6aefff",
   29314 => x"ffffff",
   29315 => x"b9d38f",
   29316 => x"3cf3cf",
   29317 => x"3cf3cf",
   29318 => x"3cf3cf",
   29319 => x"3cf3cf",
   29320 => x"3cf3cf",
   29321 => x"3cf3cf",
   29322 => x"3cf3cf",
   29323 => x"3cf3cf",
   29324 => x"3cf3cf",
   29325 => x"3cf3cf",
   29326 => x"3cf3cf",
   29327 => x"3cf3cf",
   29328 => x"3cf3cf",
   29329 => x"3cf3cf",
   29330 => x"3cf3cf",
   29331 => x"3cf3cf",
   29332 => x"3cf3cf",
   29333 => x"3cf3cf",
   29334 => x"3cf3cf",
   29335 => x"3cf3cf",
   29336 => x"3cf3ce",
   29337 => x"25afff",
   29338 => x"ffffff",
   29339 => x"ffffff",
   29340 => x"ffffff",
   29341 => x"ffffff",
   29342 => x"ffffff",
   29343 => x"ffffff",
   29344 => x"ffffff",
   29345 => x"ffffff",
   29346 => x"ffffff",
   29347 => x"ffffff",
   29348 => x"ffffff",
   29349 => x"fffa95",
   29350 => x"abffff",
   29351 => x"ffffff",
   29352 => x"ffffff",
   29353 => x"ffffff",
   29354 => x"ffffff",
   29355 => x"ffffff",
   29356 => x"ffffff",
   29357 => x"ffffff",
   29358 => x"ffffff",
   29359 => x"ffffff",
   29360 => x"ffffff",
   29361 => x"fffeb0",
   29362 => x"c30c30",
   29363 => x"c30c30",
   29364 => x"c30c30",
   29365 => x"c30c30",
   29366 => x"c30c30",
   29367 => x"c30c30",
   29368 => x"c30c30",
   29369 => x"c30c30",
   29370 => x"c30c30",
   29371 => x"c30c30",
   29372 => x"c30c30",
   29373 => x"820820",
   29374 => x"820820",
   29375 => x"820820",
   29376 => x"820820",
   29377 => x"820820",
   29378 => x"820820",
   29379 => x"820820",
   29380 => x"820820",
   29381 => x"820820",
   29382 => x"820820",
   29383 => x"820820",
   29384 => x"820820",
   29385 => x"820820",
   29386 => x"820820",
   29387 => x"820820",
   29388 => x"820820",
   29389 => x"820820",
   29390 => x"820820",
   29391 => x"820820",
   29392 => x"820820",
   29393 => x"820820",
   29394 => x"820820",
   29395 => x"820410",
   29396 => x"410410",
   29397 => x"410410",
   29398 => x"410410",
   29399 => x"410410",
   29400 => x"410410",
   29401 => x"410410",
   29402 => x"410410",
   29403 => x"410410",
   29404 => x"410410",
   29405 => x"410410",
   29406 => x"410410",
   29407 => x"410410",
   29408 => x"410410",
   29409 => x"410410",
   29410 => x"410410",
   29411 => x"410410",
   29412 => x"410410",
   29413 => x"410410",
   29414 => x"410410",
   29415 => x"410410",
   29416 => x"410410",
   29417 => x"410410",
   29418 => x"410000",
   29419 => x"000000",
   29420 => x"000000",
   29421 => x"000000",
   29422 => x"000000",
   29423 => x"000000",
   29424 => x"000000",
   29425 => x"000000",
   29426 => x"000000",
   29427 => x"000000",
   29428 => x"000000",
   29429 => x"00057f",
   29430 => x"ffffff",
   29431 => x"ffffff",
   29432 => x"ffffff",
   29433 => x"ffffff",
   29434 => x"ffffff",
   29435 => x"ffffff",
   29436 => x"ffffff",
   29437 => x"ffffff",
   29438 => x"ffffff",
   29439 => x"ffffff",
   29440 => x"ffffff",
   29441 => x"ffffff",
   29442 => x"ffffff",
   29443 => x"ffffff",
   29444 => x"ffffff",
   29445 => x"ffffff",
   29446 => x"ffffff",
   29447 => x"ffffff",
   29448 => x"ffffff",
   29449 => x"ffffff",
   29450 => x"ffffff",
   29451 => x"fd70d3",
   29452 => x"9f7cf3",
   29453 => x"cf3cf3",
   29454 => x"cf3cf3",
   29455 => x"cf3cf3",
   29456 => x"cf3cf3",
   29457 => x"cf3cf3",
   29458 => x"cf3cf3",
   29459 => x"cf3cf3",
   29460 => x"cf3cf3",
   29461 => x"cf3cf3",
   29462 => x"cf3cf3",
   29463 => x"cf3cf3",
   29464 => x"cf3cf3",
   29465 => x"cf3cf3",
   29466 => x"cf3cf3",
   29467 => x"cf3cf3",
   29468 => x"cf3cf3",
   29469 => x"cf3cf3",
   29470 => x"cf3cf3",
   29471 => x"cf3cf3",
   29472 => x"cf3cf3",
   29473 => x"deb6ae",
   29474 => x"ffffde",
   29475 => x"38f3cf",
   29476 => x"3cf3cf",
   29477 => x"3cf3cf",
   29478 => x"3cf3cf",
   29479 => x"3cf3cf",
   29480 => x"3cf3cf",
   29481 => x"3cf3cf",
   29482 => x"3cf3cf",
   29483 => x"3cf3cf",
   29484 => x"3cf3cf",
   29485 => x"3cf3cf",
   29486 => x"3cf3cf",
   29487 => x"3cf3cf",
   29488 => x"3cf3cf",
   29489 => x"3cf3cf",
   29490 => x"3cf3cf",
   29491 => x"3cf3cf",
   29492 => x"3cf3cf",
   29493 => x"3cf3cf",
   29494 => x"3cf3cf",
   29495 => x"3cf3cf",
   29496 => x"3cf286",
   29497 => x"0ebfff",
   29498 => x"ffffff",
   29499 => x"ffffff",
   29500 => x"ffffff",
   29501 => x"ffffff",
   29502 => x"ffffff",
   29503 => x"ffffff",
   29504 => x"ffffff",
   29505 => x"ffffff",
   29506 => x"ffffff",
   29507 => x"ffffff",
   29508 => x"ffffff",
   29509 => x"fffa95",
   29510 => x"abffff",
   29511 => x"ffffff",
   29512 => x"ffffff",
   29513 => x"ffffff",
   29514 => x"ffffff",
   29515 => x"ffffff",
   29516 => x"ffffff",
   29517 => x"ffffff",
   29518 => x"ffffff",
   29519 => x"ffffff",
   29520 => x"ffffff",
   29521 => x"fffeb0",
   29522 => x"c30c30",
   29523 => x"c30c30",
   29524 => x"c30c30",
   29525 => x"c30c30",
   29526 => x"c30c30",
   29527 => x"c30c30",
   29528 => x"c30c30",
   29529 => x"c30c30",
   29530 => x"c30c30",
   29531 => x"c30c30",
   29532 => x"c30c30",
   29533 => x"820820",
   29534 => x"820820",
   29535 => x"820820",
   29536 => x"820820",
   29537 => x"820820",
   29538 => x"820820",
   29539 => x"820820",
   29540 => x"820820",
   29541 => x"820820",
   29542 => x"820820",
   29543 => x"820820",
   29544 => x"820820",
   29545 => x"820820",
   29546 => x"820820",
   29547 => x"820820",
   29548 => x"820820",
   29549 => x"820820",
   29550 => x"820820",
   29551 => x"820820",
   29552 => x"820820",
   29553 => x"820820",
   29554 => x"820820",
   29555 => x"820410",
   29556 => x"410410",
   29557 => x"410410",
   29558 => x"410410",
   29559 => x"410410",
   29560 => x"410410",
   29561 => x"410410",
   29562 => x"410410",
   29563 => x"410410",
   29564 => x"410410",
   29565 => x"410410",
   29566 => x"410410",
   29567 => x"410410",
   29568 => x"410410",
   29569 => x"410410",
   29570 => x"410410",
   29571 => x"410410",
   29572 => x"410410",
   29573 => x"410410",
   29574 => x"410410",
   29575 => x"410410",
   29576 => x"410410",
   29577 => x"410410",
   29578 => x"410000",
   29579 => x"000000",
   29580 => x"000000",
   29581 => x"000000",
   29582 => x"000000",
   29583 => x"000000",
   29584 => x"000000",
   29585 => x"000000",
   29586 => x"000000",
   29587 => x"000000",
   29588 => x"000000",
   29589 => x"00057f",
   29590 => x"ffffff",
   29591 => x"ffffff",
   29592 => x"ffffff",
   29593 => x"ffffff",
   29594 => x"ffffff",
   29595 => x"ffffff",
   29596 => x"ffffff",
   29597 => x"ffffff",
   29598 => x"ffffff",
   29599 => x"ffffff",
   29600 => x"ffffff",
   29601 => x"ffffff",
   29602 => x"ffffff",
   29603 => x"ffffff",
   29604 => x"ffffff",
   29605 => x"ffffff",
   29606 => x"ffffff",
   29607 => x"ffffff",
   29608 => x"ffffff",
   29609 => x"ffffff",
   29610 => x"ffffff",
   29611 => x"fd70c3",
   29612 => x"0d79f7",
   29613 => x"cf3cf3",
   29614 => x"cf3cf3",
   29615 => x"cf3cf3",
   29616 => x"cf3cf3",
   29617 => x"cf3cf3",
   29618 => x"cf3cf3",
   29619 => x"cf3cf3",
   29620 => x"cf3cf3",
   29621 => x"cf3cf3",
   29622 => x"cf3cf3",
   29623 => x"cf3cf3",
   29624 => x"cf3cf3",
   29625 => x"cf3cf3",
   29626 => x"cf3cf3",
   29627 => x"cf3cf3",
   29628 => x"cf3cf3",
   29629 => x"cf3cf3",
   29630 => x"cf3cf3",
   29631 => x"cf3cf3",
   29632 => x"cf3cf3",
   29633 => x"cf3dd7",
   29634 => x"6ae74e",
   29635 => x"3cf3cf",
   29636 => x"3cf3cf",
   29637 => x"3cf3cf",
   29638 => x"3cf3cf",
   29639 => x"3cf3cf",
   29640 => x"3cf3cf",
   29641 => x"3cf3cf",
   29642 => x"3cf3cf",
   29643 => x"3cf3cf",
   29644 => x"3cf3cf",
   29645 => x"3cf3cf",
   29646 => x"3cf3cf",
   29647 => x"3cf3cf",
   29648 => x"3cf3cf",
   29649 => x"3cf3cf",
   29650 => x"3cf3cf",
   29651 => x"3cf3cf",
   29652 => x"3cf3cf",
   29653 => x"3cf3cf",
   29654 => x"3cf3cf",
   29655 => x"3cf3cf",
   29656 => x"38a1c3",
   29657 => x"0ebfff",
   29658 => x"ffffff",
   29659 => x"ffffff",
   29660 => x"ffffff",
   29661 => x"ffffff",
   29662 => x"ffffff",
   29663 => x"ffffff",
   29664 => x"ffffff",
   29665 => x"ffffff",
   29666 => x"ffffff",
   29667 => x"ffffff",
   29668 => x"ffffff",
   29669 => x"fffa95",
   29670 => x"abffff",
   29671 => x"ffffff",
   29672 => x"ffffff",
   29673 => x"ffffff",
   29674 => x"ffffff",
   29675 => x"ffffff",
   29676 => x"ffffff",
   29677 => x"ffffff",
   29678 => x"ffffff",
   29679 => x"ffffff",
   29680 => x"ffffff",
   29681 => x"fffeb0",
   29682 => x"c30c30",
   29683 => x"c30c30",
   29684 => x"c30c30",
   29685 => x"c30c30",
   29686 => x"c30c30",
   29687 => x"c30c30",
   29688 => x"c30c30",
   29689 => x"c30c30",
   29690 => x"c30c30",
   29691 => x"c30c30",
   29692 => x"c30c30",
   29693 => x"820820",
   29694 => x"820820",
   29695 => x"820820",
   29696 => x"820820",
   29697 => x"820820",
   29698 => x"820820",
   29699 => x"820820",
   29700 => x"820820",
   29701 => x"820820",
   29702 => x"820820",
   29703 => x"820820",
   29704 => x"820820",
   29705 => x"820820",
   29706 => x"820820",
   29707 => x"820820",
   29708 => x"820820",
   29709 => x"820820",
   29710 => x"820820",
   29711 => x"820820",
   29712 => x"820820",
   29713 => x"820820",
   29714 => x"820820",
   29715 => x"820410",
   29716 => x"410410",
   29717 => x"410410",
   29718 => x"410410",
   29719 => x"410410",
   29720 => x"410410",
   29721 => x"410410",
   29722 => x"410410",
   29723 => x"410410",
   29724 => x"410410",
   29725 => x"410410",
   29726 => x"410410",
   29727 => x"410410",
   29728 => x"410410",
   29729 => x"410410",
   29730 => x"410410",
   29731 => x"410410",
   29732 => x"410410",
   29733 => x"410410",
   29734 => x"410410",
   29735 => x"410410",
   29736 => x"410410",
   29737 => x"410410",
   29738 => x"410000",
   29739 => x"000000",
   29740 => x"000000",
   29741 => x"000000",
   29742 => x"000000",
   29743 => x"000000",
   29744 => x"000000",
   29745 => x"000000",
   29746 => x"000000",
   29747 => x"000000",
   29748 => x"000000",
   29749 => x"00057f",
   29750 => x"ffffff",
   29751 => x"ffffff",
   29752 => x"ffffff",
   29753 => x"ffffff",
   29754 => x"ffffff",
   29755 => x"ffffff",
   29756 => x"ffffff",
   29757 => x"ffffff",
   29758 => x"ffffff",
   29759 => x"ffffff",
   29760 => x"ffffff",
   29761 => x"ffffff",
   29762 => x"ffffff",
   29763 => x"ffffff",
   29764 => x"ffffff",
   29765 => x"ffffff",
   29766 => x"ffffff",
   29767 => x"ffffff",
   29768 => x"ffffff",
   29769 => x"ffffff",
   29770 => x"ffffff",
   29771 => x"fd70c3",
   29772 => x"0c30d7",
   29773 => x"af7cf3",
   29774 => x"cf3cf3",
   29775 => x"cf3cf3",
   29776 => x"cf3cf3",
   29777 => x"cf3cf3",
   29778 => x"cf3cf3",
   29779 => x"cf3cf3",
   29780 => x"cf3cf3",
   29781 => x"cf3cf3",
   29782 => x"cf3cf3",
   29783 => x"cf3cf3",
   29784 => x"cf3cf3",
   29785 => x"cf3cf3",
   29786 => x"cf3cf3",
   29787 => x"cf3cf3",
   29788 => x"cf3cf3",
   29789 => x"cf3cf3",
   29790 => x"cf3cf3",
   29791 => x"cf3cf3",
   29792 => x"cf3cf3",
   29793 => x"cf3dd7",
   29794 => x"0c624e",
   29795 => x"3cf3cf",
   29796 => x"3cf3cf",
   29797 => x"3cf3cf",
   29798 => x"3cf3cf",
   29799 => x"3cf3cf",
   29800 => x"3cf3cf",
   29801 => x"3cf3cf",
   29802 => x"3cf3cf",
   29803 => x"3cf3cf",
   29804 => x"3cf3cf",
   29805 => x"3cf3cf",
   29806 => x"3cf3cf",
   29807 => x"3cf3cf",
   29808 => x"3cf3cf",
   29809 => x"3cf3cf",
   29810 => x"3cf3cf",
   29811 => x"3cf3cf",
   29812 => x"3cf3cf",
   29813 => x"3cf3cf",
   29814 => x"3cf3cf",
   29815 => x"3cf38a",
   29816 => x"1830c3",
   29817 => x"0d7fff",
   29818 => x"ffffff",
   29819 => x"ffffff",
   29820 => x"ffffff",
   29821 => x"ffffff",
   29822 => x"ffffff",
   29823 => x"ffffff",
   29824 => x"ffffff",
   29825 => x"ffffff",
   29826 => x"ffffff",
   29827 => x"ffffff",
   29828 => x"ffffff",
   29829 => x"fffa95",
   29830 => x"abffff",
   29831 => x"ffffff",
   29832 => x"ffffff",
   29833 => x"ffffff",
   29834 => x"ffffff",
   29835 => x"ffffff",
   29836 => x"ffffff",
   29837 => x"ffffff",
   29838 => x"ffffff",
   29839 => x"ffffff",
   29840 => x"ffffff",
   29841 => x"fffeb0",
   29842 => x"c30c30",
   29843 => x"c30c30",
   29844 => x"c30c30",
   29845 => x"c30c30",
   29846 => x"c30c30",
   29847 => x"c30c30",
   29848 => x"c30c30",
   29849 => x"c30c30",
   29850 => x"c30c30",
   29851 => x"c30c30",
   29852 => x"c30c30",
   29853 => x"820820",
   29854 => x"820820",
   29855 => x"820820",
   29856 => x"820820",
   29857 => x"820820",
   29858 => x"820820",
   29859 => x"820820",
   29860 => x"820820",
   29861 => x"820820",
   29862 => x"820820",
   29863 => x"820820",
   29864 => x"820820",
   29865 => x"820820",
   29866 => x"820820",
   29867 => x"820820",
   29868 => x"820820",
   29869 => x"820820",
   29870 => x"820820",
   29871 => x"820820",
   29872 => x"820820",
   29873 => x"820820",
   29874 => x"820820",
   29875 => x"820810",
   29876 => x"410410",
   29877 => x"410410",
   29878 => x"410410",
   29879 => x"410410",
   29880 => x"410410",
   29881 => x"410410",
   29882 => x"410410",
   29883 => x"410410",
   29884 => x"410410",
   29885 => x"410410",
   29886 => x"410410",
   29887 => x"410410",
   29888 => x"410410",
   29889 => x"410410",
   29890 => x"410410",
   29891 => x"410410",
   29892 => x"410410",
   29893 => x"410410",
   29894 => x"410410",
   29895 => x"410410",
   29896 => x"410410",
   29897 => x"410410",
   29898 => x"410000",
   29899 => x"000000",
   29900 => x"000000",
   29901 => x"000000",
   29902 => x"000000",
   29903 => x"000000",
   29904 => x"000000",
   29905 => x"000000",
   29906 => x"000000",
   29907 => x"000000",
   29908 => x"000000",
   29909 => x"00057f",
   29910 => x"ffffff",
   29911 => x"ffffff",
   29912 => x"ffffff",
   29913 => x"ffffff",
   29914 => x"ffffff",
   29915 => x"ffffff",
   29916 => x"ffffff",
   29917 => x"ffffff",
   29918 => x"ffffff",
   29919 => x"ffffff",
   29920 => x"ffffff",
   29921 => x"ffffff",
   29922 => x"ffffff",
   29923 => x"ffffff",
   29924 => x"ffffff",
   29925 => x"ffffff",
   29926 => x"ffffff",
   29927 => x"ffffff",
   29928 => x"ffffff",
   29929 => x"ffffff",
   29930 => x"ffffff",
   29931 => x"ad70c3",
   29932 => x"0c30c3",
   29933 => x"0d79f7",
   29934 => x"df3cf3",
   29935 => x"cf3cf3",
   29936 => x"cf3cf3",
   29937 => x"cf3cf3",
   29938 => x"cf3cf3",
   29939 => x"cf3cf3",
   29940 => x"cf3cf3",
   29941 => x"cf3cf3",
   29942 => x"cf3cf3",
   29943 => x"cf3cf3",
   29944 => x"cf3cf3",
   29945 => x"cf3cf3",
   29946 => x"cf3cf3",
   29947 => x"cf3cf3",
   29948 => x"cf3cf3",
   29949 => x"cf3cf3",
   29950 => x"cf3cf3",
   29951 => x"cf3cf3",
   29952 => x"cf3cf7",
   29953 => x"dd70c3",
   29954 => x"0c30c7",
   29955 => x"28e3cf",
   29956 => x"3cf3cf",
   29957 => x"3cf3cf",
   29958 => x"3cf3cf",
   29959 => x"3cf3cf",
   29960 => x"3cf3cf",
   29961 => x"3cf3cf",
   29962 => x"3cf3cf",
   29963 => x"3cf3cf",
   29964 => x"3cf3cf",
   29965 => x"3cf3cf",
   29966 => x"3cf3cf",
   29967 => x"3cf3cf",
   29968 => x"3cf3cf",
   29969 => x"3cf3cf",
   29970 => x"3cf3cf",
   29971 => x"3cf3cf",
   29972 => x"3cf3cf",
   29973 => x"3cf3cf",
   29974 => x"3cf3cf",
   29975 => x"38a1c3",
   29976 => x"0c30c3",
   29977 => x"0d7fff",
   29978 => x"ffffff",
   29979 => x"ffffff",
   29980 => x"ffffff",
   29981 => x"ffffff",
   29982 => x"ffffff",
   29983 => x"ffffff",
   29984 => x"ffffff",
   29985 => x"ffffff",
   29986 => x"ffffff",
   29987 => x"ffffff",
   29988 => x"ffffff",
   29989 => x"fffa95",
   29990 => x"abffff",
   29991 => x"ffffff",
   29992 => x"ffffff",
   29993 => x"ffffff",
   29994 => x"ffffff",
   29995 => x"ffffff",
   29996 => x"ffffff",
   29997 => x"ffffff",
   29998 => x"ffffff",
   29999 => x"ffffff",
   30000 => x"ffffff",
   30001 => x"fffeb5",
   30002 => x"c30c30",
   30003 => x"c30c30",
   30004 => x"c30c30",
   30005 => x"c30c30",
   30006 => x"c30c30",
   30007 => x"c30c30",
   30008 => x"c30c30",
   30009 => x"c30c30",
   30010 => x"c30c30",
   30011 => x"c30c30",
   30012 => x"c30c30",
   30013 => x"c30c30",
   30014 => x"c30c20",
   30015 => x"820820",
   30016 => x"820820",
   30017 => x"820820",
   30018 => x"820820",
   30019 => x"820820",
   30020 => x"820820",
   30021 => x"820820",
   30022 => x"820820",
   30023 => x"820820",
   30024 => x"820820",
   30025 => x"820820",
   30026 => x"820820",
   30027 => x"820820",
   30028 => x"820820",
   30029 => x"820820",
   30030 => x"820820",
   30031 => x"820820",
   30032 => x"820820",
   30033 => x"820820",
   30034 => x"820820",
   30035 => x"820820",
   30036 => x"820820",
   30037 => x"820820",
   30038 => x"820820",
   30039 => x"820820",
   30040 => x"820820",
   30041 => x"410410",
   30042 => x"410410",
   30043 => x"410410",
   30044 => x"410410",
   30045 => x"410410",
   30046 => x"410410",
   30047 => x"410410",
   30048 => x"410410",
   30049 => x"410410",
   30050 => x"410410",
   30051 => x"410410",
   30052 => x"410410",
   30053 => x"410410",
   30054 => x"410410",
   30055 => x"410410",
   30056 => x"410410",
   30057 => x"410410",
   30058 => x"410410",
   30059 => x"410410",
   30060 => x"410410",
   30061 => x"410410",
   30062 => x"410410",
   30063 => x"410410",
   30064 => x"410410",
   30065 => x"410410",
   30066 => x"410410",
   30067 => x"400000",
   30068 => x"000000",
   30069 => x"000abf",
   30070 => x"ffffff",
   30071 => x"ffffff",
   30072 => x"ffffff",
   30073 => x"ffffff",
   30074 => x"ffffff",
   30075 => x"ffffff",
   30076 => x"ffffff",
   30077 => x"ffffff",
   30078 => x"ffffff",
   30079 => x"ffffff",
   30080 => x"ffffff",
   30081 => x"ffffff",
   30082 => x"ffffff",
   30083 => x"ffffff",
   30084 => x"ffffff",
   30085 => x"ffffff",
   30086 => x"ffffff",
   30087 => x"ffffff",
   30088 => x"ffffff",
   30089 => x"ffffff",
   30090 => x"ffffff",
   30091 => x"ad70c3",
   30092 => x"0c30c3",
   30093 => x"0c30d3",
   30094 => x"5fbdf3",
   30095 => x"cf3cf3",
   30096 => x"cf3cf3",
   30097 => x"cf3cf3",
   30098 => x"cf3cf3",
   30099 => x"cf3cf3",
   30100 => x"cf3cf3",
   30101 => x"cf3cf3",
   30102 => x"cf3cf3",
   30103 => x"cf3cf3",
   30104 => x"cf3cf3",
   30105 => x"cf3cf3",
   30106 => x"cf3cf3",
   30107 => x"cf3cf3",
   30108 => x"cf3cf3",
   30109 => x"cf3cf3",
   30110 => x"cf3cf3",
   30111 => x"cf3cf3",
   30112 => x"cf79d7",
   30113 => x"0c30c3",
   30114 => x"0c30c3",
   30115 => x"0c728e",
   30116 => x"3cf3cf",
   30117 => x"3cf3cf",
   30118 => x"3cf3cf",
   30119 => x"3cf3cf",
   30120 => x"3cf3cf",
   30121 => x"3cf3cf",
   30122 => x"3cf3cf",
   30123 => x"3cf3cf",
   30124 => x"3cf3cf",
   30125 => x"3cf3cf",
   30126 => x"3cf3cf",
   30127 => x"3cf3cf",
   30128 => x"3cf3cf",
   30129 => x"3cf3cf",
   30130 => x"3cf3cf",
   30131 => x"3cf3cf",
   30132 => x"3cf3cf",
   30133 => x"3cf3cf",
   30134 => x"3ce38a",
   30135 => x"1c30c3",
   30136 => x"0c30c3",
   30137 => x"0d7fff",
   30138 => x"ffffff",
   30139 => x"ffffff",
   30140 => x"ffffff",
   30141 => x"ffffff",
   30142 => x"ffffff",
   30143 => x"ffffff",
   30144 => x"ffffff",
   30145 => x"ffffff",
   30146 => x"ffffff",
   30147 => x"ffffff",
   30148 => x"ffffff",
   30149 => x"fffa95",
   30150 => x"abffff",
   30151 => x"ffffff",
   30152 => x"ffffff",
   30153 => x"ffffff",
   30154 => x"ffffff",
   30155 => x"ffffff",
   30156 => x"ffffff",
   30157 => x"ffffff",
   30158 => x"ffffff",
   30159 => x"ffffff",
   30160 => x"ffffff",
   30161 => x"ffffff",
   30162 => x"ffffff",
   30163 => x"ffffff",
   30164 => x"ffffff",
   30165 => x"ffffff",
   30166 => x"ffffff",
   30167 => x"ffffff",
   30168 => x"ffffff",
   30169 => x"ffffff",
   30170 => x"ffffff",
   30171 => x"ffffff",
   30172 => x"ffffff",
   30173 => x"ffffff",
   30174 => x"ffffff",
   30175 => x"ffffff",
   30176 => x"ffffff",
   30177 => x"ffffff",
   30178 => x"ffffff",
   30179 => x"ffffff",
   30180 => x"ffffff",
   30181 => x"ffffff",
   30182 => x"ffffff",
   30183 => x"ffffff",
   30184 => x"ffffff",
   30185 => x"ffffff",
   30186 => x"ffffff",
   30187 => x"ffffff",
   30188 => x"ffffff",
   30189 => x"ffffff",
   30190 => x"ffffff",
   30191 => x"ffffff",
   30192 => x"ffffff",
   30193 => x"ffffff",
   30194 => x"ffffff",
   30195 => x"ffffff",
   30196 => x"ffffff",
   30197 => x"ffffff",
   30198 => x"ffffff",
   30199 => x"ffffff",
   30200 => x"ffffff",
   30201 => x"ffffff",
   30202 => x"ffffff",
   30203 => x"ffffff",
   30204 => x"ffffff",
   30205 => x"ffffff",
   30206 => x"ffffff",
   30207 => x"ffffff",
   30208 => x"ffffff",
   30209 => x"ffffff",
   30210 => x"ffffff",
   30211 => x"ffffff",
   30212 => x"ffffff",
   30213 => x"ffffff",
   30214 => x"ffffff",
   30215 => x"ffffff",
   30216 => x"ffffff",
   30217 => x"ffffff",
   30218 => x"ffffff",
   30219 => x"ffffff",
   30220 => x"ffffff",
   30221 => x"ffffff",
   30222 => x"ffffff",
   30223 => x"ffffff",
   30224 => x"ffffff",
   30225 => x"ffffff",
   30226 => x"ffffff",
   30227 => x"ffffff",
   30228 => x"ffffff",
   30229 => x"ffffff",
   30230 => x"ffffff",
   30231 => x"ffffff",
   30232 => x"ffffff",
   30233 => x"ffffff",
   30234 => x"ffffff",
   30235 => x"ffffff",
   30236 => x"ffffff",
   30237 => x"ffffff",
   30238 => x"ffffff",
   30239 => x"ffffff",
   30240 => x"ffffff",
   30241 => x"ffffff",
   30242 => x"ffffff",
   30243 => x"ffffff",
   30244 => x"ffffff",
   30245 => x"ffffff",
   30246 => x"ffffff",
   30247 => x"ffffff",
   30248 => x"ffffff",
   30249 => x"ffffff",
   30250 => x"ffffff",
   30251 => x"ad70c3",
   30252 => x"0c30c3",
   30253 => x"0c30c3",
   30254 => x"0d35eb",
   30255 => x"df7cf3",
   30256 => x"cf3cf3",
   30257 => x"cf3cf3",
   30258 => x"cf3cf3",
   30259 => x"cf3cf3",
   30260 => x"cf3cf3",
   30261 => x"cf3cf3",
   30262 => x"cf3cf3",
   30263 => x"cf3cf3",
   30264 => x"cf3cf3",
   30265 => x"cf3cf3",
   30266 => x"cf3cf3",
   30267 => x"cf3cf3",
   30268 => x"cf3cf3",
   30269 => x"cf3cf3",
   30270 => x"cf3cf3",
   30271 => x"cf3de7",
   30272 => x"5d30c3",
   30273 => x"0c30c3",
   30274 => x"0c30c3",
   30275 => x"0c30c7",
   30276 => x"28e38f",
   30277 => x"3cf3cf",
   30278 => x"3cf3cf",
   30279 => x"3cf3cf",
   30280 => x"3cf3cf",
   30281 => x"3cf3cf",
   30282 => x"3cf3cf",
   30283 => x"3cf3cf",
   30284 => x"3cf3cf",
   30285 => x"3cf3cf",
   30286 => x"3cf3cf",
   30287 => x"3cf3cf",
   30288 => x"3cf3cf",
   30289 => x"3cf3cf",
   30290 => x"3cf3cf",
   30291 => x"3cf3cf",
   30292 => x"3cf3cf",
   30293 => x"3cf3ce",
   30294 => x"2461c3",
   30295 => x"0c30c3",
   30296 => x"0c30c3",
   30297 => x"0d7fff",
   30298 => x"ffffff",
   30299 => x"ffffff",
   30300 => x"ffffff",
   30301 => x"ffffff",
   30302 => x"ffffff",
   30303 => x"ffffff",
   30304 => x"ffffff",
   30305 => x"ffffff",
   30306 => x"ffffff",
   30307 => x"ffffff",
   30308 => x"ffffff",
   30309 => x"fffa95",
   30310 => x"abffff",
   30311 => x"ffffff",
   30312 => x"ffffff",
   30313 => x"ffffff",
   30314 => x"ffffff",
   30315 => x"ffffff",
   30316 => x"ffffff",
   30317 => x"ffffff",
   30318 => x"ffffff",
   30319 => x"ffffff",
   30320 => x"ffffff",
   30321 => x"ffffff",
   30322 => x"ffffff",
   30323 => x"ffffff",
   30324 => x"ffffff",
   30325 => x"ffffff",
   30326 => x"ffffff",
   30327 => x"ffffff",
   30328 => x"ffffff",
   30329 => x"ffffff",
   30330 => x"ffffff",
   30331 => x"ffffff",
   30332 => x"ffffff",
   30333 => x"ffffff",
   30334 => x"ffffff",
   30335 => x"ffffff",
   30336 => x"ffffff",
   30337 => x"ffffff",
   30338 => x"ffffff",
   30339 => x"ffffff",
   30340 => x"ffffff",
   30341 => x"ffffff",
   30342 => x"ffffff",
   30343 => x"ffffff",
   30344 => x"ffffff",
   30345 => x"ffffff",
   30346 => x"ffffff",
   30347 => x"ffffff",
   30348 => x"ffffff",
   30349 => x"ffffff",
   30350 => x"ffffff",
   30351 => x"ffffff",
   30352 => x"ffffff",
   30353 => x"ffffff",
   30354 => x"ffffff",
   30355 => x"ffffff",
   30356 => x"ffffff",
   30357 => x"ffffff",
   30358 => x"ffffff",
   30359 => x"ffffff",
   30360 => x"ffffff",
   30361 => x"ffffff",
   30362 => x"ffffff",
   30363 => x"ffffff",
   30364 => x"ffffff",
   30365 => x"ffffff",
   30366 => x"ffffff",
   30367 => x"ffffff",
   30368 => x"ffffff",
   30369 => x"ffffff",
   30370 => x"ffffff",
   30371 => x"ffffff",
   30372 => x"ffffff",
   30373 => x"ffffff",
   30374 => x"ffffff",
   30375 => x"ffffff",
   30376 => x"ffffff",
   30377 => x"ffffff",
   30378 => x"ffffff",
   30379 => x"ffffff",
   30380 => x"ffffff",
   30381 => x"ffffff",
   30382 => x"ffffff",
   30383 => x"ffffff",
   30384 => x"ffffff",
   30385 => x"ffffff",
   30386 => x"ffffff",
   30387 => x"ffffff",
   30388 => x"ffffff",
   30389 => x"ffffff",
   30390 => x"ffffff",
   30391 => x"ffffff",
   30392 => x"ffffff",
   30393 => x"ffffff",
   30394 => x"ffffff",
   30395 => x"ffffff",
   30396 => x"ffffff",
   30397 => x"ffffff",
   30398 => x"ffffff",
   30399 => x"ffffff",
   30400 => x"ffffff",
   30401 => x"ffffff",
   30402 => x"ffffff",
   30403 => x"ffffff",
   30404 => x"ffffff",
   30405 => x"ffffff",
   30406 => x"ffffff",
   30407 => x"ffffff",
   30408 => x"ffffff",
   30409 => x"ffffff",
   30410 => x"ffffff",
   30411 => x"ac30c3",
   30412 => x"0c30c3",
   30413 => x"0c30c3",
   30414 => x"0c30c3",
   30415 => x"5e7df7",
   30416 => x"cf3cf3",
   30417 => x"cf3cf3",
   30418 => x"cf3cf3",
   30419 => x"cf3cf3",
   30420 => x"cf3cf3",
   30421 => x"cf3cf3",
   30422 => x"cf3cf3",
   30423 => x"cf3cf3",
   30424 => x"cf3cf3",
   30425 => x"cf3cf3",
   30426 => x"cf3cf3",
   30427 => x"cf3cf3",
   30428 => x"cf3cf3",
   30429 => x"cf3cf3",
   30430 => x"cf3cf7",
   30431 => x"de75d3",
   30432 => x"0c30c3",
   30433 => x"0c30c3",
   30434 => x"0c30c3",
   30435 => x"0c30c3",
   30436 => x"0c718a",
   30437 => x"38e3cf",
   30438 => x"3cf3cf",
   30439 => x"3cf3cf",
   30440 => x"3cf3cf",
   30441 => x"3cf3cf",
   30442 => x"3cf3cf",
   30443 => x"3cf3cf",
   30444 => x"3cf3cf",
   30445 => x"3cf3cf",
   30446 => x"3cf3cf",
   30447 => x"3cf3cf",
   30448 => x"3cf3cf",
   30449 => x"3cf3cf",
   30450 => x"3cf3cf",
   30451 => x"3cf3cf",
   30452 => x"3cf3cf",
   30453 => x"38e286",
   30454 => x"1c30c3",
   30455 => x"0c30c3",
   30456 => x"0c30c3",
   30457 => x"0d7fff",
   30458 => x"ffffff",
   30459 => x"ffffff",
   30460 => x"ffffff",
   30461 => x"ffffff",
   30462 => x"ffffff",
   30463 => x"ffffff",
   30464 => x"ffffff",
   30465 => x"ffffff",
   30466 => x"ffffff",
   30467 => x"ffffff",
   30468 => x"ffffff",
   30469 => x"fffa95",
   30470 => x"abffff",
   30471 => x"ffffff",
   30472 => x"ffffff",
   30473 => x"ffffff",
   30474 => x"ffffff",
   30475 => x"ffffff",
   30476 => x"ffffff",
   30477 => x"ffffff",
   30478 => x"ffffff",
   30479 => x"ffffff",
   30480 => x"ffffff",
   30481 => x"ffffff",
   30482 => x"ffffff",
   30483 => x"ffffff",
   30484 => x"ffffff",
   30485 => x"ffffff",
   30486 => x"ffffff",
   30487 => x"ffffff",
   30488 => x"ffffff",
   30489 => x"ffffff",
   30490 => x"ffffff",
   30491 => x"ffffff",
   30492 => x"ffffff",
   30493 => x"ffffff",
   30494 => x"ffffff",
   30495 => x"ffffff",
   30496 => x"ffffff",
   30497 => x"ffffff",
   30498 => x"ffffff",
   30499 => x"ffffff",
   30500 => x"ffffff",
   30501 => x"ffffff",
   30502 => x"ffffff",
   30503 => x"ffffff",
   30504 => x"ffffff",
   30505 => x"ffffff",
   30506 => x"ffffff",
   30507 => x"ffffff",
   30508 => x"ffffff",
   30509 => x"ffffff",
   30510 => x"ffffff",
   30511 => x"ffffff",
   30512 => x"ffffff",
   30513 => x"ffffff",
   30514 => x"ffffff",
   30515 => x"ffffff",
   30516 => x"ffffff",
   30517 => x"ffffff",
   30518 => x"ffffff",
   30519 => x"ffffff",
   30520 => x"ffffff",
   30521 => x"ffffff",
   30522 => x"ffffff",
   30523 => x"ffffff",
   30524 => x"ffffff",
   30525 => x"ffffff",
   30526 => x"ffffff",
   30527 => x"ffffff",
   30528 => x"ffffff",
   30529 => x"ffffff",
   30530 => x"ffffff",
   30531 => x"ffffff",
   30532 => x"ffffff",
   30533 => x"ffffff",
   30534 => x"ffffff",
   30535 => x"ffffff",
   30536 => x"ffffff",
   30537 => x"ffffff",
   30538 => x"ffffff",
   30539 => x"ffffff",
   30540 => x"ffffff",
   30541 => x"ffffff",
   30542 => x"ffffff",
   30543 => x"ffffff",
   30544 => x"ffffff",
   30545 => x"ffffff",
   30546 => x"ffffff",
   30547 => x"ffffff",
   30548 => x"ffffff",
   30549 => x"ffffff",
   30550 => x"ffffff",
   30551 => x"ffffff",
   30552 => x"ffffff",
   30553 => x"ffffff",
   30554 => x"ffffff",
   30555 => x"ffffff",
   30556 => x"ffffff",
   30557 => x"ffffff",
   30558 => x"ffffff",
   30559 => x"ffffff",
   30560 => x"ffffff",
   30561 => x"ffffff",
   30562 => x"ffffff",
   30563 => x"ffffff",
   30564 => x"ffffff",
   30565 => x"ffffff",
   30566 => x"ffffff",
   30567 => x"ffffff",
   30568 => x"ffffff",
   30569 => x"ffffff",
   30570 => x"ffffff",
   30571 => x"ac30c3",
   30572 => x"0c30c3",
   30573 => x"0c30c3",
   30574 => x"0c30c3",
   30575 => x"0c35d7",
   30576 => x"9f7df3",
   30577 => x"cf3cf3",
   30578 => x"cf3cf3",
   30579 => x"cf3cf3",
   30580 => x"cf3cf3",
   30581 => x"cf3cf3",
   30582 => x"cf3cf3",
   30583 => x"cf3cf3",
   30584 => x"cf3cf3",
   30585 => x"cf3cf3",
   30586 => x"cf3cf3",
   30587 => x"cf3cf3",
   30588 => x"cf3cf3",
   30589 => x"cf3cf3",
   30590 => x"df79d7",
   30591 => x"4c30c3",
   30592 => x"0c30c3",
   30593 => x"0c30c3",
   30594 => x"0c30c3",
   30595 => x"0c30c3",
   30596 => x"0c30c3",
   30597 => x"1c628e",
   30598 => x"38f3cf",
   30599 => x"3cf3cf",
   30600 => x"3cf3cf",
   30601 => x"3cf3cf",
   30602 => x"3cf3cf",
   30603 => x"3cf3cf",
   30604 => x"3cf3cf",
   30605 => x"3cf3cf",
   30606 => x"3cf3cf",
   30607 => x"3cf3cf",
   30608 => x"3cf3cf",
   30609 => x"3cf3cf",
   30610 => x"3cf3cf",
   30611 => x"3cf3cf",
   30612 => x"3ce38a",
   30613 => x"1860c3",
   30614 => x"0c30c3",
   30615 => x"0c30c3",
   30616 => x"0c30c3",
   30617 => x"0d7fff",
   30618 => x"ffffff",
   30619 => x"ffffff",
   30620 => x"ffffff",
   30621 => x"ffffff",
   30622 => x"ffffff",
   30623 => x"ffffff",
   30624 => x"ffffff",
   30625 => x"ffffff",
   30626 => x"ffffff",
   30627 => x"ffffff",
   30628 => x"ffffff",
   30629 => x"fffa95",
   30630 => x"abffff",
   30631 => x"ffffff",
   30632 => x"ffffff",
   30633 => x"ffffff",
   30634 => x"ffffff",
   30635 => x"ffffff",
   30636 => x"ffffff",
   30637 => x"ffffff",
   30638 => x"ffffff",
   30639 => x"ffffff",
   30640 => x"ffffff",
   30641 => x"ffffff",
   30642 => x"ffffff",
   30643 => x"ffffff",
   30644 => x"ffffff",
   30645 => x"ffffff",
   30646 => x"ffffff",
   30647 => x"ffffff",
   30648 => x"ffffff",
   30649 => x"ffffff",
   30650 => x"ffffff",
   30651 => x"ffffff",
   30652 => x"ffffff",
   30653 => x"ffffff",
   30654 => x"ffffff",
   30655 => x"ffffff",
   30656 => x"ffffff",
   30657 => x"ffffff",
   30658 => x"ffffff",
   30659 => x"ffffff",
   30660 => x"ffffff",
   30661 => x"ffffff",
   30662 => x"ffffff",
   30663 => x"ffffff",
   30664 => x"ffffff",
   30665 => x"ffffff",
   30666 => x"ffffff",
   30667 => x"ffffff",
   30668 => x"ffffff",
   30669 => x"ffffff",
   30670 => x"ffffff",
   30671 => x"ffffff",
   30672 => x"ffffff",
   30673 => x"ffffff",
   30674 => x"ffffff",
   30675 => x"ffffff",
   30676 => x"ffffff",
   30677 => x"ffffff",
   30678 => x"ffffff",
   30679 => x"ffffff",
   30680 => x"ffffff",
   30681 => x"ffffff",
   30682 => x"ffffff",
   30683 => x"ffffff",
   30684 => x"ffffff",
   30685 => x"ffffff",
   30686 => x"ffffff",
   30687 => x"ffffff",
   30688 => x"ffffff",
   30689 => x"ffffff",
   30690 => x"ffffff",
   30691 => x"ffffff",
   30692 => x"ffffff",
   30693 => x"ffffff",
   30694 => x"ffffff",
   30695 => x"ffffff",
   30696 => x"ffffff",
   30697 => x"ffffff",
   30698 => x"ffffff",
   30699 => x"ffffff",
   30700 => x"ffffff",
   30701 => x"ffffff",
   30702 => x"ffffff",
   30703 => x"ffffff",
   30704 => x"ffffff",
   30705 => x"ffffff",
   30706 => x"ffffff",
   30707 => x"ffffff",
   30708 => x"ffffff",
   30709 => x"ffffff",
   30710 => x"ffffff",
   30711 => x"ffffff",
   30712 => x"ffffff",
   30713 => x"ffffff",
   30714 => x"ffffff",
   30715 => x"ffffff",
   30716 => x"ffffff",
   30717 => x"ffffff",
   30718 => x"ffffff",
   30719 => x"ffffff",
   30720 => x"ffffff",
   30721 => x"ffffff",
   30722 => x"ffffff",
   30723 => x"ffffff",
   30724 => x"ffffff",
   30725 => x"ffffff",
   30726 => x"ffffff",
   30727 => x"ffffff",
   30728 => x"ffffff",
   30729 => x"ffffff",
   30730 => x"ffffff",
   30731 => x"ac30c3",
   30732 => x"0c30c3",
   30733 => x"0c30c3",
   30734 => x"0c30c3",
   30735 => x"0c30c3",
   30736 => x"0d35e7",
   30737 => x"9f7df3",
   30738 => x"cf3cf3",
   30739 => x"cf3cf3",
   30740 => x"cf3cf3",
   30741 => x"cf3cf3",
   30742 => x"cf3cf3",
   30743 => x"cf3cf3",
   30744 => x"cf3cf3",
   30745 => x"cf3cf3",
   30746 => x"cf3cf3",
   30747 => x"cf3cf3",
   30748 => x"cf3cf3",
   30749 => x"df79e7",
   30750 => x"5d70c3",
   30751 => x"0c30c3",
   30752 => x"0c30c3",
   30753 => x"0c30c3",
   30754 => x"0c30c3",
   30755 => x"0c30c3",
   30756 => x"0c30c3",
   30757 => x"0c30c6",
   30758 => x"18a38e",
   30759 => x"3cf3cf",
   30760 => x"3cf3cf",
   30761 => x"3cf3cf",
   30762 => x"3cf3cf",
   30763 => x"3cf3cf",
   30764 => x"3cf3cf",
   30765 => x"3cf3cf",
   30766 => x"3cf3cf",
   30767 => x"3cf3cf",
   30768 => x"3cf3cf",
   30769 => x"3cf3cf",
   30770 => x"3cf3cf",
   30771 => x"3ce38e",
   30772 => x"286183",
   30773 => x"0c30c3",
   30774 => x"0c30c3",
   30775 => x"0c30c3",
   30776 => x"0c30c3",
   30777 => x"0d7fff",
   30778 => x"ffffff",
   30779 => x"ffffff",
   30780 => x"ffffff",
   30781 => x"ffffff",
   30782 => x"ffffff",
   30783 => x"ffffff",
   30784 => x"ffffff",
   30785 => x"ffffff",
   30786 => x"ffffff",
   30787 => x"ffffff",
   30788 => x"ffffff",
   30789 => x"fffa95",
   30790 => x"abffff",
   30791 => x"ffffff",
   30792 => x"ffffff",
   30793 => x"ffffff",
   30794 => x"ffffff",
   30795 => x"ffffff",
   30796 => x"ffffff",
   30797 => x"ffffff",
   30798 => x"ffffff",
   30799 => x"ffffff",
   30800 => x"ffffff",
   30801 => x"ffffff",
   30802 => x"ffffff",
   30803 => x"ffffff",
   30804 => x"ffffff",
   30805 => x"ffffff",
   30806 => x"ffffff",
   30807 => x"ffffff",
   30808 => x"ffffff",
   30809 => x"ffffff",
   30810 => x"ffffff",
   30811 => x"ffffff",
   30812 => x"ffffff",
   30813 => x"ffffff",
   30814 => x"ffffff",
   30815 => x"ffffff",
   30816 => x"ffffff",
   30817 => x"ffffff",
   30818 => x"ffffff",
   30819 => x"ffffff",
   30820 => x"ffffff",
   30821 => x"ffffff",
   30822 => x"ffffff",
   30823 => x"ffffff",
   30824 => x"ffffff",
   30825 => x"ffffff",
   30826 => x"ffffff",
   30827 => x"ffffff",
   30828 => x"ffffff",
   30829 => x"ffffff",
   30830 => x"ffffff",
   30831 => x"ffffff",
   30832 => x"ffffff",
   30833 => x"ffffff",
   30834 => x"ffffff",
   30835 => x"ffffff",
   30836 => x"ffffff",
   30837 => x"ffffff",
   30838 => x"ffffff",
   30839 => x"ffffff",
   30840 => x"ffffff",
   30841 => x"ffffff",
   30842 => x"ffffff",
   30843 => x"ffffff",
   30844 => x"ffffff",
   30845 => x"ffffff",
   30846 => x"ffffff",
   30847 => x"ffffff",
   30848 => x"ffffff",
   30849 => x"ffffff",
   30850 => x"ffffff",
   30851 => x"ffffff",
   30852 => x"ffffff",
   30853 => x"ffffff",
   30854 => x"ffffff",
   30855 => x"ffffff",
   30856 => x"ffffff",
   30857 => x"ffffff",
   30858 => x"ffffff",
   30859 => x"ffffff",
   30860 => x"ffffff",
   30861 => x"ffffff",
   30862 => x"ffffff",
   30863 => x"ffffff",
   30864 => x"ffffff",
   30865 => x"ffffff",
   30866 => x"ffffff",
   30867 => x"ffffff",
   30868 => x"ffffff",
   30869 => x"ffffff",
   30870 => x"ffffff",
   30871 => x"ffffff",
   30872 => x"ffffff",
   30873 => x"ffffff",
   30874 => x"ffffff",
   30875 => x"ffffff",
   30876 => x"ffffff",
   30877 => x"ffffff",
   30878 => x"ffffff",
   30879 => x"ffffff",
   30880 => x"ffffff",
   30881 => x"ffffff",
   30882 => x"ffffff",
   30883 => x"ffffff",
   30884 => x"ffffff",
   30885 => x"ffffff",
   30886 => x"ffffff",
   30887 => x"ffffff",
   30888 => x"ffffff",
   30889 => x"ffffff",
   30890 => x"ffffff",
   30891 => x"ad70c3",
   30892 => x"0c30c3",
   30893 => x"0c30c3",
   30894 => x"0c30c3",
   30895 => x"0c30c3",
   30896 => x"0c30c3",
   30897 => x"5d75e7",
   30898 => x"9f7df3",
   30899 => x"cf3cf3",
   30900 => x"cf3cf3",
   30901 => x"cf3cf3",
   30902 => x"cf3cf3",
   30903 => x"cf3cf3",
   30904 => x"cf3cf3",
   30905 => x"cf3cf3",
   30906 => x"cf3cf3",
   30907 => x"cf3cf3",
   30908 => x"df79e7",
   30909 => x"5d75c3",
   30910 => x"0c30c3",
   30911 => x"0c30c3",
   30912 => x"0c30c3",
   30913 => x"0c30c3",
   30914 => x"0c30c3",
   30915 => x"0c30c3",
   30916 => x"0c30c3",
   30917 => x"0c30c3",
   30918 => x"0c6186",
   30919 => x"28a38e",
   30920 => x"3cf3cf",
   30921 => x"3cf3cf",
   30922 => x"3cf3cf",
   30923 => x"3cf3cf",
   30924 => x"3cf3cf",
   30925 => x"3cf3cf",
   30926 => x"3cf3cf",
   30927 => x"3cf3cf",
   30928 => x"3cf3cf",
   30929 => x"3cf3cf",
   30930 => x"3ce38e",
   30931 => x"28a186",
   30932 => x"1830c3",
   30933 => x"0c30c3",
   30934 => x"0c30c3",
   30935 => x"0c30c3",
   30936 => x"0c30c3",
   30937 => x"0d7fff",
   30938 => x"ffffff",
   30939 => x"ffffff",
   30940 => x"ffffff",
   30941 => x"ffffff",
   30942 => x"ffffff",
   30943 => x"ffffff",
   30944 => x"ffffff",
   30945 => x"ffffff",
   30946 => x"ffffff",
   30947 => x"ffffff",
   30948 => x"ffffff",
   30949 => x"fffa95",
   30950 => x"abffff",
   30951 => x"ffffff",
   30952 => x"ffffff",
   30953 => x"ffffff",
   30954 => x"ffffff",
   30955 => x"ffffff",
   30956 => x"ffffff",
   30957 => x"ffffff",
   30958 => x"ffffff",
   30959 => x"ffffff",
   30960 => x"ffffff",
   30961 => x"ffffff",
   30962 => x"ffffff",
   30963 => x"ffffff",
   30964 => x"ffffff",
   30965 => x"ffffff",
   30966 => x"ffffff",
   30967 => x"ffffff",
   30968 => x"ffffff",
   30969 => x"ffffff",
   30970 => x"ffffff",
   30971 => x"ffffff",
   30972 => x"ffffff",
   30973 => x"ffffff",
   30974 => x"ffffff",
   30975 => x"ffffff",
   30976 => x"ffffff",
   30977 => x"ffffff",
   30978 => x"ffffff",
   30979 => x"ffffff",
   30980 => x"ffffff",
   30981 => x"ffffff",
   30982 => x"ffffff",
   30983 => x"ffffff",
   30984 => x"ffffff",
   30985 => x"ffffff",
   30986 => x"ffffff",
   30987 => x"ffffff",
   30988 => x"ffffff",
   30989 => x"ffffff",
   30990 => x"ffffff",
   30991 => x"ffffff",
   30992 => x"ffffff",
   30993 => x"ffffff",
   30994 => x"ffffff",
   30995 => x"ffffff",
   30996 => x"ffffff",
   30997 => x"ffffff",
   30998 => x"ffffff",
   30999 => x"ffffff",
   31000 => x"ffffff",
   31001 => x"ffffff",
   31002 => x"ffffff",
   31003 => x"ffffff",
   31004 => x"ffffff",
   31005 => x"ffffff",
   31006 => x"ffffff",
   31007 => x"ffffff",
   31008 => x"ffffff",
   31009 => x"ffffff",
   31010 => x"ffffff",
   31011 => x"ffffff",
   31012 => x"ffffff",
   31013 => x"ffffff",
   31014 => x"ffffff",
   31015 => x"ffffff",
   31016 => x"ffffff",
   31017 => x"ffffff",
   31018 => x"ffffff",
   31019 => x"ffffff",
   31020 => x"ffffff",
   31021 => x"ffffff",
   31022 => x"ffffff",
   31023 => x"ffffff",
   31024 => x"ffffff",
   31025 => x"ffffff",
   31026 => x"ffffff",
   31027 => x"ffffff",
   31028 => x"ffffff",
   31029 => x"ffffff",
   31030 => x"ffffff",
   31031 => x"ffffff",
   31032 => x"ffffff",
   31033 => x"ffffff",
   31034 => x"ffffff",
   31035 => x"ffffff",
   31036 => x"ffffff",
   31037 => x"ffffff",
   31038 => x"ffffff",
   31039 => x"ffffff",
   31040 => x"ffffff",
   31041 => x"ffffff",
   31042 => x"ffffff",
   31043 => x"ffffff",
   31044 => x"ffffff",
   31045 => x"ffffff",
   31046 => x"ffffff",
   31047 => x"ffffff",
   31048 => x"ffffff",
   31049 => x"ffffff",
   31050 => x"ffffff",
   31051 => x"ad70c3",
   31052 => x"0c30c3",
   31053 => x"0c30c3",
   31054 => x"0c30c3",
   31055 => x"0c30c3",
   31056 => x"0c30c3",
   31057 => x"0c30c3",
   31058 => x"5d75e7",
   31059 => x"9f7df7",
   31060 => x"df3cf3",
   31061 => x"cf3cf3",
   31062 => x"cf3cf3",
   31063 => x"cf3cf3",
   31064 => x"cf3cf3",
   31065 => x"cf3cf3",
   31066 => x"df7df7",
   31067 => x"df79e7",
   31068 => x"5d75c3",
   31069 => x"0c30c3",
   31070 => x"0c30c3",
   31071 => x"0c30c3",
   31072 => x"0c30c3",
   31073 => x"0c30c3",
   31074 => x"0c30c3",
   31075 => x"0c30c3",
   31076 => x"0c30c3",
   31077 => x"0c30c3",
   31078 => x"0c30c3",
   31079 => x"0c6186",
   31080 => x"28a38e",
   31081 => x"38f3cf",
   31082 => x"3cf3cf",
   31083 => x"3cf3cf",
   31084 => x"3cf3cf",
   31085 => x"3cf3cf",
   31086 => x"3cf3cf",
   31087 => x"3cf3cf",
   31088 => x"3cf3ce",
   31089 => x"38e38e",
   31090 => x"28a186",
   31091 => x"1830c3",
   31092 => x"0c30c3",
   31093 => x"0c30c3",
   31094 => x"0c30c3",
   31095 => x"0c30c3",
   31096 => x"0c30c3",
   31097 => x"0d7fff",
   31098 => x"ffffff",
   31099 => x"ffffff",
   31100 => x"ffffff",
   31101 => x"ffffff",
   31102 => x"ffffff",
   31103 => x"ffffff",
   31104 => x"ffffff",
   31105 => x"ffffff",
   31106 => x"ffffff",
   31107 => x"ffffff",
   31108 => x"ffffff",
   31109 => x"fffa95",
   31110 => x"abffff",
   31111 => x"ffffff",
   31112 => x"ffffff",
   31113 => x"ffffff",
   31114 => x"ffffff",
   31115 => x"ffffff",
   31116 => x"ffffff",
   31117 => x"ffffff",
   31118 => x"ffffff",
   31119 => x"ffffff",
   31120 => x"ffffff",
   31121 => x"ffffff",
   31122 => x"ffffff",
   31123 => x"ffffff",
   31124 => x"ffffff",
   31125 => x"ffffff",
   31126 => x"ffffff",
   31127 => x"ffffff",
   31128 => x"ffffff",
   31129 => x"ffffff",
   31130 => x"ffffff",
   31131 => x"ffffff",
   31132 => x"ffffff",
   31133 => x"ffffff",
   31134 => x"ffffff",
   31135 => x"ffffff",
   31136 => x"ffffff",
   31137 => x"ffffff",
   31138 => x"ffffff",
   31139 => x"ffffff",
   31140 => x"ffffff",
   31141 => x"ffffff",
   31142 => x"ffffff",
   31143 => x"ffffff",
   31144 => x"ffffff",
   31145 => x"ffffff",
   31146 => x"ffffff",
   31147 => x"ffffff",
   31148 => x"ffffff",
   31149 => x"ffffff",
   31150 => x"ffffff",
   31151 => x"ffffff",
   31152 => x"ffffff",
   31153 => x"ffffff",
   31154 => x"ffffff",
   31155 => x"ffffff",
   31156 => x"ffffff",
   31157 => x"ffffff",
   31158 => x"ffffff",
   31159 => x"ffffff",
   31160 => x"ffffff",
   31161 => x"ffffff",
   31162 => x"ffffff",
   31163 => x"ffffff",
   31164 => x"ffffff",
   31165 => x"ffffff",
   31166 => x"ffffff",
   31167 => x"ffffff",
   31168 => x"ffffff",
   31169 => x"ffffff",
   31170 => x"ffffff",
   31171 => x"ffffff",
   31172 => x"ffffff",
   31173 => x"ffffff",
   31174 => x"ffffff",
   31175 => x"ffffff",
   31176 => x"ffffff",
   31177 => x"ffffff",
   31178 => x"ffffff",
   31179 => x"ffffff",
   31180 => x"ffffff",
   31181 => x"ffffff",
   31182 => x"ffffff",
   31183 => x"ffffff",
   31184 => x"ffffff",
   31185 => x"ffffff",
   31186 => x"ffffff",
   31187 => x"ffffff",
   31188 => x"ffffff",
   31189 => x"ffffff",
   31190 => x"ffffff",
   31191 => x"ffffff",
   31192 => x"ffffff",
   31193 => x"ffffff",
   31194 => x"ffffff",
   31195 => x"ffffff",
   31196 => x"ffffff",
   31197 => x"ffffff",
   31198 => x"ffffff",
   31199 => x"ffffff",
   31200 => x"ffffff",
   31201 => x"ffffff",
   31202 => x"ffffff",
   31203 => x"ffffff",
   31204 => x"ffffff",
   31205 => x"ffffff",
   31206 => x"ffffff",
   31207 => x"ffffff",
   31208 => x"ffffff",
   31209 => x"ffffff",
   31210 => x"ffffff",
   31211 => x"ad70c3",
   31212 => x"0c30c3",
   31213 => x"0c30c3",
   31214 => x"0c30c3",
   31215 => x"0c30c3",
   31216 => x"0c30c3",
   31217 => x"0c30c3",
   31218 => x"0c30c3",
   31219 => x"5d75d7",
   31220 => x"9e79e7",
   31221 => x"df7df7",
   31222 => x"df7df7",
   31223 => x"df7df7",
   31224 => x"df7df7",
   31225 => x"9e79e7",
   31226 => x"9e75d7",
   31227 => x"5d75c3",
   31228 => x"0c30c3",
   31229 => x"0c30c3",
   31230 => x"0c30c3",
   31231 => x"0c30c3",
   31232 => x"0c30c3",
   31233 => x"0c30c3",
   31234 => x"0c30c3",
   31235 => x"0c30c3",
   31236 => x"0c30c3",
   31237 => x"0c30c3",
   31238 => x"0c30c3",
   31239 => x"0c30c3",
   31240 => x"0c6186",
   31241 => x"18a28a",
   31242 => x"38e38e",
   31243 => x"3cf3cf",
   31244 => x"3cf3cf",
   31245 => x"3cf3cf",
   31246 => x"3cf3ce",
   31247 => x"38e38e",
   31248 => x"38e28a",
   31249 => x"286186",
   31250 => x"1830c3",
   31251 => x"0c30c3",
   31252 => x"0c30c3",
   31253 => x"0c30c3",
   31254 => x"0c30c3",
   31255 => x"0c30c3",
   31256 => x"0c30c3",
   31257 => x"0d7fff",
   31258 => x"ffffff",
   31259 => x"ffffff",
   31260 => x"ffffff",
   31261 => x"ffffff",
   31262 => x"ffffff",
   31263 => x"ffffff",
   31264 => x"ffffff",
   31265 => x"ffffff",
   31266 => x"ffffff",
   31267 => x"ffffff",
   31268 => x"ffffff",
   31269 => x"fffa95",
   31270 => x"abffff",
   31271 => x"ffffff",
   31272 => x"ffffff",
   31273 => x"ffffff",
   31274 => x"ffffff",
   31275 => x"ffffff",
   31276 => x"ffffff",
   31277 => x"ffffff",
   31278 => x"ffffff",
   31279 => x"ffffff",
   31280 => x"ffffff",
   31281 => x"ffffff",
   31282 => x"ffffff",
   31283 => x"ffffff",
   31284 => x"ffffff",
   31285 => x"ffffff",
   31286 => x"ffffff",
   31287 => x"ffffff",
   31288 => x"ffffff",
   31289 => x"ffffff",
   31290 => x"ffffff",
   31291 => x"ffffff",
   31292 => x"ffffff",
   31293 => x"ffffff",
   31294 => x"ffffff",
   31295 => x"ffffff",
   31296 => x"ffffff",
   31297 => x"ffffff",
   31298 => x"ffffff",
   31299 => x"ffffff",
   31300 => x"ffffff",
   31301 => x"ffffff",
   31302 => x"ffffff",
   31303 => x"ffffff",
   31304 => x"ffffff",
   31305 => x"ffffff",
   31306 => x"ffffff",
   31307 => x"ffffff",
   31308 => x"ffffff",
   31309 => x"ffffff",
   31310 => x"ffffff",
   31311 => x"ffffff",
   31312 => x"ffffff",
   31313 => x"ffffff",
   31314 => x"ffffff",
   31315 => x"ffffff",
   31316 => x"ffffff",
   31317 => x"ffffff",
   31318 => x"ffffff",
   31319 => x"ffffff",
   31320 => x"ffffff",
   31321 => x"ffffff",
   31322 => x"ffffff",
   31323 => x"ffffff",
   31324 => x"ffffff",
   31325 => x"ffffff",
   31326 => x"ffffff",
   31327 => x"ffffff",
   31328 => x"ffffff",
   31329 => x"ffffff",
   31330 => x"ffffff",
   31331 => x"ffffff",
   31332 => x"ffffff",
   31333 => x"ffffff",
   31334 => x"ffffff",
   31335 => x"ffffff",
   31336 => x"ffffff",
   31337 => x"ffffff",
   31338 => x"ffffff",
   31339 => x"ffffff",
   31340 => x"ffffff",
   31341 => x"ffffff",
   31342 => x"ffffff",
   31343 => x"ffffff",
   31344 => x"ffffff",
   31345 => x"ffffff",
   31346 => x"ffffff",
   31347 => x"ffffff",
   31348 => x"ffffff",
   31349 => x"ffffff",
   31350 => x"ffffff",
   31351 => x"ffffff",
   31352 => x"ffffff",
   31353 => x"ffffff",
   31354 => x"ffffff",
   31355 => x"ffffff",
   31356 => x"ffffff",
   31357 => x"ffffff",
   31358 => x"ffffff",
   31359 => x"ffffff",
   31360 => x"ffffff",
   31361 => x"ffffff",
   31362 => x"ffffff",
   31363 => x"ffffff",
   31364 => x"ffffff",
   31365 => x"ffffff",
   31366 => x"ffffff",
   31367 => x"ffffff",
   31368 => x"ffffff",
   31369 => x"ffffff",
   31370 => x"ffffff",
   31371 => x"ad70c3",
   31372 => x"0c30c3",
   31373 => x"0c30c3",
   31374 => x"0c30c3",
   31375 => x"0c30c3",
   31376 => x"0c30c3",
   31377 => x"0c30c3",
   31378 => x"0c30c3",
   31379 => x"0c30c3",
   31380 => x"0c35d7",
   31381 => x"5d75d7",
   31382 => x"5d75d7",
   31383 => x"5d75d7",
   31384 => x"5d75d7",
   31385 => x"5d75c3",
   31386 => x"0c30c3",
   31387 => x"0c30c3",
   31388 => x"0c30c3",
   31389 => x"0c30c3",
   31390 => x"0c30c3",
   31391 => x"0c30c3",
   31392 => x"0c30c3",
   31393 => x"0c30c3",
   31394 => x"0c30c3",
   31395 => x"0c30c3",
   31396 => x"0c30c3",
   31397 => x"0c30c3",
   31398 => x"0c30c3",
   31399 => x"0c30c3",
   31400 => x"0c30c3",
   31401 => x"0c3186",
   31402 => x"18618a",
   31403 => x"28a28a",
   31404 => x"28a28a",
   31405 => x"28a28a",
   31406 => x"28a28a",
   31407 => x"28a286",
   31408 => x"186182",
   31409 => x"0c30c3",
   31410 => x"0c30c3",
   31411 => x"0c30c3",
   31412 => x"0c30c3",
   31413 => x"0c30c3",
   31414 => x"0c30c3",
   31415 => x"0c30c3",
   31416 => x"0c30c3",
   31417 => x"0d7fff",
   31418 => x"ffffff",
   31419 => x"ffffff",
   31420 => x"ffffff",
   31421 => x"ffffff",
   31422 => x"ffffff",
   31423 => x"ffffff",
   31424 => x"ffffff",
   31425 => x"ffffff",
   31426 => x"ffffff",
   31427 => x"ffffff",
   31428 => x"ffffff",
   31429 => x"fffa95",
   31430 => x"abffff",
   31431 => x"ffffff",
   31432 => x"ffffff",
   31433 => x"ffffff",
   31434 => x"ffffff",
   31435 => x"ffffff",
   31436 => x"ffffff",
   31437 => x"ffffff",
   31438 => x"ffffff",
   31439 => x"ffffff",
   31440 => x"ffffff",
   31441 => x"ffffff",
   31442 => x"ffffff",
   31443 => x"ffffff",
   31444 => x"ffffff",
   31445 => x"ffffff",
   31446 => x"ffffff",
   31447 => x"ffffff",
   31448 => x"ffffff",
   31449 => x"ffffff",
   31450 => x"ffffff",
   31451 => x"ffffff",
   31452 => x"ffffff",
   31453 => x"ffffff",
   31454 => x"ffffff",
   31455 => x"ffffff",
   31456 => x"ffffff",
   31457 => x"ffffff",
   31458 => x"ffffff",
   31459 => x"ffffff",
   31460 => x"ffffff",
   31461 => x"ffffff",
   31462 => x"ffffff",
   31463 => x"ffffff",
   31464 => x"ffffff",
   31465 => x"ffffff",
   31466 => x"ffffff",
   31467 => x"ffffff",
   31468 => x"ffffff",
   31469 => x"ffffff",
   31470 => x"ffffff",
   31471 => x"ffffff",
   31472 => x"ffffff",
   31473 => x"ffffff",
   31474 => x"ffffff",
   31475 => x"ffffff",
   31476 => x"ffffff",
   31477 => x"ffffff",
   31478 => x"ffffff",
   31479 => x"ffffff",
   31480 => x"ffffff",
   31481 => x"ffffff",
   31482 => x"ffffff",
   31483 => x"ffffff",
   31484 => x"ffffff",
   31485 => x"ffffff",
   31486 => x"ffffff",
   31487 => x"ffffff",
   31488 => x"ffffff",
   31489 => x"ffffff",
   31490 => x"ffffff",
   31491 => x"ffffff",
   31492 => x"ffffff",
   31493 => x"ffffff",
   31494 => x"ffffff",
   31495 => x"ffffff",
   31496 => x"ffffff",
   31497 => x"ffffff",
   31498 => x"ffffff",
   31499 => x"ffffff",
   31500 => x"ffffff",
   31501 => x"ffffff",
   31502 => x"ffffff",
   31503 => x"ffffff",
   31504 => x"ffffff",
   31505 => x"ffffff",
   31506 => x"ffffff",
   31507 => x"ffffff",
   31508 => x"ffffff",
   31509 => x"ffffff",
   31510 => x"ffffff",
   31511 => x"ffffff",
   31512 => x"ffffff",
   31513 => x"ffffff",
   31514 => x"ffffff",
   31515 => x"ffffff",
   31516 => x"ffffff",
   31517 => x"ffffff",
   31518 => x"ffffff",
   31519 => x"ffffff",
   31520 => x"ffffff",
   31521 => x"ffffff",
   31522 => x"ffffff",
   31523 => x"ffffff",
   31524 => x"ffffff",
   31525 => x"ffffff",
   31526 => x"ffffff",
   31527 => x"ffffff",
   31528 => x"ffffff",
   31529 => x"ffffff",
   31530 => x"ffffff",
   31531 => x"fd70c3",
   31532 => x"0c30c3",
   31533 => x"0c30c3",
   31534 => x"0c30c3",
   31535 => x"0c30c3",
   31536 => x"0c30c3",
   31537 => x"0c30c3",
   31538 => x"0c30c3",
   31539 => x"0c30c3",
   31540 => x"0c30c3",
   31541 => x"0c30c3",
   31542 => x"0c30c3",
   31543 => x"0c30c3",
   31544 => x"0c30c3",
   31545 => x"0c30c3",
   31546 => x"0c30c3",
   31547 => x"0c30c3",
   31548 => x"0c30c3",
   31549 => x"0c30c3",
   31550 => x"0c30c3",
   31551 => x"0c30c3",
   31552 => x"0c30c3",
   31553 => x"0c30c3",
   31554 => x"0c30c3",
   31555 => x"0c30c3",
   31556 => x"0c30c3",
   31557 => x"0c30c3",
   31558 => x"0c30c3",
   31559 => x"0c30c3",
   31560 => x"0c30c3",
   31561 => x"0c30c3",
   31562 => x"0c30c3",
   31563 => x"0c30c3",
   31564 => x"086186",
   31565 => x"186186",
   31566 => x"1820c3",
   31567 => x"0c30c3",
   31568 => x"0c30c3",
   31569 => x"0c30c3",
   31570 => x"0c30c3",
   31571 => x"0c30c3",
   31572 => x"0c30c3",
   31573 => x"0c30c3",
   31574 => x"0c30c3",
   31575 => x"0c30c3",
   31576 => x"0c30c3",
   31577 => x"0d7fff",
   31578 => x"ffffff",
   31579 => x"ffffff",
   31580 => x"ffffff",
   31581 => x"ffffff",
   31582 => x"ffffff",
   31583 => x"ffffff",
   31584 => x"ffffff",
   31585 => x"ffffff",
   31586 => x"ffffff",
   31587 => x"ffffff",
   31588 => x"ffffff",
   31589 => x"fffa95",
   31590 => x"abffff",
   31591 => x"ffffff",
   31592 => x"ffffff",
   31593 => x"ffffff",
   31594 => x"ffffff",
   31595 => x"ffffff",
   31596 => x"ffffff",
   31597 => x"ffffff",
   31598 => x"ffffff",
   31599 => x"ffffff",
   31600 => x"ffffff",
   31601 => x"ffffff",
   31602 => x"ffffff",
   31603 => x"ffffff",
   31604 => x"ffffff",
   31605 => x"ffffff",
   31606 => x"ffffff",
   31607 => x"ffffff",
   31608 => x"ffffff",
   31609 => x"ffffff",
   31610 => x"ffffff",
   31611 => x"ffffff",
   31612 => x"ffffff",
   31613 => x"ffffff",
   31614 => x"ffffff",
   31615 => x"ffffff",
   31616 => x"ffffff",
   31617 => x"ffffff",
   31618 => x"ffffff",
   31619 => x"ffffff",
   31620 => x"ffffff",
   31621 => x"ffffff",
   31622 => x"ffffff",
   31623 => x"ffffff",
   31624 => x"ffffff",
   31625 => x"ffffff",
   31626 => x"ffffff",
   31627 => x"ffffff",
   31628 => x"ffffff",
   31629 => x"ffffff",
   31630 => x"ffffff",
   31631 => x"ffffff",
   31632 => x"ffffff",
   31633 => x"ffffff",
   31634 => x"ffffff",
   31635 => x"ffffff",
   31636 => x"ffffff",
   31637 => x"ffffff",
   31638 => x"ffffff",
   31639 => x"ffffff",
   31640 => x"ffffff",
   31641 => x"ffffff",
   31642 => x"ffffff",
   31643 => x"ffffff",
   31644 => x"ffffff",
   31645 => x"ffffff",
   31646 => x"ffffff",
   31647 => x"ffffff",
   31648 => x"ffffff",
   31649 => x"ffffff",
   31650 => x"ffffff",
   31651 => x"ffffff",
   31652 => x"ffffff",
   31653 => x"ffffff",
   31654 => x"ffffff",
   31655 => x"ffffff",
   31656 => x"ffffff",
   31657 => x"ffffff",
   31658 => x"ffffff",
   31659 => x"ffffff",
   31660 => x"ffffff",
   31661 => x"ffffff",
   31662 => x"ffffff",
   31663 => x"ffffff",
   31664 => x"ffffff",
   31665 => x"ffffff",
   31666 => x"ffffff",
   31667 => x"ffffff",
   31668 => x"ffffff",
   31669 => x"ffffff",
   31670 => x"ffffff",
   31671 => x"ffffff",
   31672 => x"ffffff",
   31673 => x"ffffff",
   31674 => x"ffffff",
   31675 => x"ffffff",
   31676 => x"ffffff",
   31677 => x"ffffff",
   31678 => x"ffffff",
   31679 => x"ffffff",
   31680 => x"ffffff",
   31681 => x"ffffff",
   31682 => x"ffffff",
   31683 => x"ffffff",
   31684 => x"ffffff",
   31685 => x"ffffff",
   31686 => x"ffffff",
   31687 => x"ffffff",
   31688 => x"ffffff",
   31689 => x"ffffff",
   31690 => x"ffffff",
   31691 => x"fd70c3",
   31692 => x"0c30c3",
   31693 => x"0c30c3",
   31694 => x"0c30c3",
   31695 => x"0c30c3",
   31696 => x"0c30c3",
   31697 => x"0c30c3",
   31698 => x"0c30c3",
   31699 => x"0c30c3",
   31700 => x"0c30c3",
   31701 => x"0c30c3",
   31702 => x"0c30c3",
   31703 => x"0c30c3",
   31704 => x"0c30c3",
   31705 => x"0c30c3",
   31706 => x"0c30c3",
   31707 => x"0c30c3",
   31708 => x"0c30c3",
   31709 => x"0c30c3",
   31710 => x"0c30c3",
   31711 => x"0c30c3",
   31712 => x"0c30c3",
   31713 => x"0c30c3",
   31714 => x"0c30c3",
   31715 => x"0c30c3",
   31716 => x"0c30c3",
   31717 => x"0c30c3",
   31718 => x"0c30c3",
   31719 => x"0c30c3",
   31720 => x"0c30c3",
   31721 => x"0c30c3",
   31722 => x"0c30c3",
   31723 => x"0c30c3",
   31724 => x"0c30c3",
   31725 => x"0c30c3",
   31726 => x"0c30c3",
   31727 => x"0c30c3",
   31728 => x"0c30c3",
   31729 => x"0c30c3",
   31730 => x"0c30c3",
   31731 => x"0c30c3",
   31732 => x"0c30c3",
   31733 => x"0c30c3",
   31734 => x"0c30c3",
   31735 => x"0c30c3",
   31736 => x"0c30c3",
   31737 => x"0ebfff",
   31738 => x"ffffff",
   31739 => x"ffffff",
   31740 => x"ffffff",
   31741 => x"ffffff",
   31742 => x"ffffff",
   31743 => x"ffffff",
   31744 => x"ffffff",
   31745 => x"ffffff",
   31746 => x"ffffff",
   31747 => x"ffffff",
   31748 => x"ffffff",
   31749 => x"fffa95",
   31750 => x"abffff",
   31751 => x"ffffff",
   31752 => x"ffffff",
   31753 => x"ffffff",
   31754 => x"ffffff",
   31755 => x"ffffff",
   31756 => x"ffffff",
   31757 => x"ffffff",
   31758 => x"ffffff",
   31759 => x"ffffff",
   31760 => x"ffffff",
   31761 => x"ffffff",
   31762 => x"ffffff",
   31763 => x"ffffff",
   31764 => x"ffffff",
   31765 => x"ffffff",
   31766 => x"ffffff",
   31767 => x"ffffff",
   31768 => x"ffffff",
   31769 => x"ffffff",
   31770 => x"ffffff",
   31771 => x"ffffff",
   31772 => x"ffffff",
   31773 => x"ffffff",
   31774 => x"ffffff",
   31775 => x"ffffff",
   31776 => x"ffffff",
   31777 => x"ffffff",
   31778 => x"ffffff",
   31779 => x"ffffff",
   31780 => x"ffffff",
   31781 => x"ffffff",
   31782 => x"ffffff",
   31783 => x"ffffff",
   31784 => x"ffffff",
   31785 => x"ffffff",
   31786 => x"ffffff",
   31787 => x"ffffff",
   31788 => x"ffffff",
   31789 => x"ffffff",
   31790 => x"ffffff",
   31791 => x"ffffff",
   31792 => x"ffffff",
   31793 => x"ffffff",
   31794 => x"ffffff",
   31795 => x"ffffff",
   31796 => x"ffffff",
   31797 => x"ffffff",
   31798 => x"ffffff",
   31799 => x"ffffff",
   31800 => x"ffffff",
   31801 => x"ffffff",
   31802 => x"ffffff",
   31803 => x"ffffff",
   31804 => x"ffffff",
   31805 => x"ffffff",
   31806 => x"ffffff",
   31807 => x"ffffff",
   31808 => x"ffffff",
   31809 => x"ffffff",
   31810 => x"ffffff",
   31811 => x"ffffff",
   31812 => x"ffffff",
   31813 => x"ffffff",
   31814 => x"ffffff",
   31815 => x"ffffff",
   31816 => x"ffffff",
   31817 => x"ffffff",
   31818 => x"ffffff",
   31819 => x"ffffff",
   31820 => x"ffffff",
   31821 => x"ffffff",
   31822 => x"ffffff",
   31823 => x"ffffff",
   31824 => x"ffffff",
   31825 => x"ffffff",
   31826 => x"ffffff",
   31827 => x"ffffff",
   31828 => x"ffffff",
   31829 => x"ffffff",
   31830 => x"ffffff",
   31831 => x"ffffff",
   31832 => x"ffffff",
   31833 => x"ffffff",
   31834 => x"ffffff",
   31835 => x"ffffff",
   31836 => x"ffffff",
   31837 => x"ffffff",
   31838 => x"ffffff",
   31839 => x"ffffff",
   31840 => x"ffffff",
   31841 => x"ffffff",
   31842 => x"ffffff",
   31843 => x"ffffff",
   31844 => x"ffffff",
   31845 => x"ffffff",
   31846 => x"ffffff",
   31847 => x"ffffff",
   31848 => x"ffffff",
   31849 => x"ffffff",
   31850 => x"ffffff",
   31851 => x"fd70c3",
   31852 => x"0c30c3",
   31853 => x"0c30c3",
   31854 => x"0c30c3",
   31855 => x"0c30c3",
   31856 => x"0c30c3",
   31857 => x"0c30c3",
   31858 => x"0c30c3",
   31859 => x"0c30c3",
   31860 => x"0c30c3",
   31861 => x"0c30c3",
   31862 => x"0c30c3",
   31863 => x"0c30c3",
   31864 => x"0c30c3",
   31865 => x"0c30c3",
   31866 => x"0c30c3",
   31867 => x"0c30c3",
   31868 => x"0c30c3",
   31869 => x"0c30c3",
   31870 => x"0c30c3",
   31871 => x"0c30c3",
   31872 => x"0c30c3",
   31873 => x"0c30c3",
   31874 => x"0c30c3",
   31875 => x"0c30c3",
   31876 => x"0c30c3",
   31877 => x"0c30c3",
   31878 => x"0c30c3",
   31879 => x"0c30c3",
   31880 => x"0c30c3",
   31881 => x"0c30c3",
   31882 => x"0c30c3",
   31883 => x"0c30c3",
   31884 => x"0c30c3",
   31885 => x"0c30c3",
   31886 => x"0c30c3",
   31887 => x"0c30c3",
   31888 => x"0c30c3",
   31889 => x"0c30c3",
   31890 => x"0c30c3",
   31891 => x"0c30c3",
   31892 => x"0c30c3",
   31893 => x"0c30c3",
   31894 => x"0c30c3",
   31895 => x"0c30c3",
   31896 => x"0c30c3",
   31897 => x"0ebfff",
   31898 => x"ffffff",
   31899 => x"ffffff",
   31900 => x"ffffff",
   31901 => x"ffffff",
   31902 => x"ffffff",
   31903 => x"ffffff",
   31904 => x"ffffff",
   31905 => x"ffffff",
   31906 => x"ffffff",
   31907 => x"ffffff",
   31908 => x"ffffff",
   31909 => x"fffa95",
   31910 => x"abffff",
   31911 => x"ffffff",
   31912 => x"ffffff",
   31913 => x"ffffff",
   31914 => x"ffffff",
   31915 => x"ffffff",
   31916 => x"ffffff",
   31917 => x"ffffff",
   31918 => x"ffffff",
   31919 => x"ffffff",
   31920 => x"ffffff",
   31921 => x"ffffff",
   31922 => x"ffffff",
   31923 => x"ffffff",
   31924 => x"ffffff",
   31925 => x"ffffff",
   31926 => x"ffffff",
   31927 => x"ffffff",
   31928 => x"ffffff",
   31929 => x"ffffff",
   31930 => x"ffffff",
   31931 => x"ffffff",
   31932 => x"ffffff",
   31933 => x"ffffff",
   31934 => x"ffffff",
   31935 => x"ffffff",
   31936 => x"ffffff",
   31937 => x"ffffff",
   31938 => x"ffffff",
   31939 => x"ffffff",
   31940 => x"ffffff",
   31941 => x"ffffff",
   31942 => x"ffffff",
   31943 => x"ffffff",
   31944 => x"ffffff",
   31945 => x"ffffff",
   31946 => x"ffffff",
   31947 => x"ffffff",
   31948 => x"ffffff",
   31949 => x"ffffff",
   31950 => x"ffffff",
   31951 => x"ffffff",
   31952 => x"ffffff",
   31953 => x"ffffff",
   31954 => x"ffffff",
   31955 => x"ffffff",
   31956 => x"ffffff",
   31957 => x"ffffff",
   31958 => x"ffffff",
   31959 => x"ffffff",
   31960 => x"ffffff",
   31961 => x"ffffff",
   31962 => x"ffffff",
   31963 => x"ffffff",
   31964 => x"ffffff",
   31965 => x"ffffff",
   31966 => x"ffffff",
   31967 => x"ffffff",
   31968 => x"ffffff",
   31969 => x"ffffff",
   31970 => x"ffffff",
   31971 => x"ffffff",
   31972 => x"ffffff",
   31973 => x"ffffff",
   31974 => x"ffffff",
   31975 => x"ffffff",
   31976 => x"ffffff",
   31977 => x"ffffff",
   31978 => x"ffffff",
   31979 => x"ffffff",
   31980 => x"ffffff",
   31981 => x"ffffff",
   31982 => x"ffffff",
   31983 => x"ffffff",
   31984 => x"ffffff",
   31985 => x"ffffff",
   31986 => x"ffffff",
   31987 => x"ffffff",
   31988 => x"ffffff",
   31989 => x"ffffff",
   31990 => x"ffffff",
   31991 => x"ffffff",
   31992 => x"ffffff",
   31993 => x"ffffff",
   31994 => x"ffffff",
   31995 => x"ffffff",
   31996 => x"ffffff",
   31997 => x"ffffff",
   31998 => x"ffffff",
   31999 => x"ffffff",
   32000 => x"ffffff",
   32001 => x"ffffff",
   32002 => x"ffffff",
   32003 => x"ffffff",
   32004 => x"ffffff",
   32005 => x"ffffff",
   32006 => x"ffffff",
   32007 => x"ffffff",
   32008 => x"ffffff",
   32009 => x"ffffff",
   32010 => x"ffffff",
   32011 => x"fd70c3",
   32012 => x"0c30c3",
   32013 => x"0c30c3",
   32014 => x"0c30c3",
   32015 => x"0c30c3",
   32016 => x"0c30c3",
   32017 => x"0c30c3",
   32018 => x"0c30c3",
   32019 => x"0c30c3",
   32020 => x"0c30c3",
   32021 => x"0c30c3",
   32022 => x"0c30c3",
   32023 => x"0c30c3",
   32024 => x"0c30c3",
   32025 => x"0c30c3",
   32026 => x"0c30c3",
   32027 => x"0c30c3",
   32028 => x"0c30c3",
   32029 => x"0c30c3",
   32030 => x"0c30c3",
   32031 => x"0c30c3",
   32032 => x"0c30c3",
   32033 => x"0c30c3",
   32034 => x"0c30c3",
   32035 => x"0c30c3",
   32036 => x"0c30c3",
   32037 => x"0c30c3",
   32038 => x"0c30c3",
   32039 => x"0c30c3",
   32040 => x"0c30c3",
   32041 => x"0c30c3",
   32042 => x"0c30c3",
   32043 => x"0c30c3",
   32044 => x"0c30c3",
   32045 => x"0c30c3",
   32046 => x"0c30c3",
   32047 => x"0c30c3",
   32048 => x"0c30c3",
   32049 => x"0c30c3",
   32050 => x"0c30c3",
   32051 => x"0c30c3",
   32052 => x"0c30c3",
   32053 => x"0c30c3",
   32054 => x"0c30c3",
   32055 => x"0c30c3",
   32056 => x"0c30c3",
   32057 => x"0ebfff",
   32058 => x"ffffff",
   32059 => x"ffffff",
   32060 => x"ffffff",
   32061 => x"ffffff",
   32062 => x"ffffff",
   32063 => x"ffffff",
   32064 => x"ffffff",
   32065 => x"ffffff",
   32066 => x"ffffff",
   32067 => x"ffffff",
   32068 => x"ffffff",
   32069 => x"fffa95",
   32070 => x"abffff",
   32071 => x"ffffff",
   32072 => x"ffffff",
   32073 => x"ffffff",
   32074 => x"ffffff",
   32075 => x"ffffff",
   32076 => x"ffffff",
   32077 => x"ffffff",
   32078 => x"ffffff",
   32079 => x"ffffff",
   32080 => x"ffffff",
   32081 => x"ffffff",
   32082 => x"ffffff",
   32083 => x"ffffff",
   32084 => x"ffffff",
   32085 => x"ffffff",
   32086 => x"ffffff",
   32087 => x"ffffff",
   32088 => x"ffffff",
   32089 => x"ffffff",
   32090 => x"ffffff",
   32091 => x"ffffff",
   32092 => x"ffffff",
   32093 => x"ffffff",
   32094 => x"ffffff",
   32095 => x"ffffff",
   32096 => x"ffffff",
   32097 => x"ffffff",
   32098 => x"ffffff",
   32099 => x"ffffff",
   32100 => x"ffffff",
   32101 => x"ffffff",
   32102 => x"ffffff",
   32103 => x"ffffff",
   32104 => x"ffffff",
   32105 => x"ffffff",
   32106 => x"ffffff",
   32107 => x"ffffff",
   32108 => x"ffffff",
   32109 => x"ffffff",
   32110 => x"ffffff",
   32111 => x"ffffff",
   32112 => x"ffffff",
   32113 => x"ffffff",
   32114 => x"ffffff",
   32115 => x"ffffff",
   32116 => x"ffffff",
   32117 => x"ffffff",
   32118 => x"ffffff",
   32119 => x"ffffff",
   32120 => x"ffffff",
   32121 => x"ffffff",
   32122 => x"ffffff",
   32123 => x"ffffff",
   32124 => x"ffffff",
   32125 => x"ffffff",
   32126 => x"ffffff",
   32127 => x"ffffff",
   32128 => x"ffffff",
   32129 => x"ffffff",
   32130 => x"ffffff",
   32131 => x"ffffff",
   32132 => x"ffffff",
   32133 => x"ffffff",
   32134 => x"ffffff",
   32135 => x"ffffff",
   32136 => x"ffffff",
   32137 => x"ffffff",
   32138 => x"ffffff",
   32139 => x"ffffff",
   32140 => x"ffffff",
   32141 => x"ffffff",
   32142 => x"ffffff",
   32143 => x"ffffff",
   32144 => x"ffffff",
   32145 => x"ffffff",
   32146 => x"ffffff",
   32147 => x"ffffff",
   32148 => x"ffffff",
   32149 => x"ffffff",
   32150 => x"ffffff",
   32151 => x"ffffff",
   32152 => x"ffffff",
   32153 => x"ffffff",
   32154 => x"ffffff",
   32155 => x"ffffff",
   32156 => x"ffffff",
   32157 => x"ffffff",
   32158 => x"ffffff",
   32159 => x"ffffff",
   32160 => x"ffffff",
   32161 => x"ffffff",
   32162 => x"ffffff",
   32163 => x"ffffff",
   32164 => x"ffffff",
   32165 => x"ffffff",
   32166 => x"ffffff",
   32167 => x"ffffff",
   32168 => x"ffffff",
   32169 => x"ffffff",
   32170 => x"ffffff",
   32171 => x"fd70c3",
   32172 => x"0c30c3",
   32173 => x"0c30c3",
   32174 => x"0c30c3",
   32175 => x"0c30c3",
   32176 => x"0c30c3",
   32177 => x"0c30c3",
   32178 => x"0c30c3",
   32179 => x"0c30c3",
   32180 => x"0c30c3",
   32181 => x"0c30c3",
   32182 => x"0c30c3",
   32183 => x"0c30c3",
   32184 => x"0c30c3",
   32185 => x"0c30c3",
   32186 => x"0c30c3",
   32187 => x"0c30c3",
   32188 => x"0c30c3",
   32189 => x"0c30c3",
   32190 => x"0c30c3",
   32191 => x"0c30c3",
   32192 => x"0c30c3",
   32193 => x"0c30c3",
   32194 => x"0c30c3",
   32195 => x"0c30c3",
   32196 => x"0c30c3",
   32197 => x"0c30c3",
   32198 => x"0c30c3",
   32199 => x"0c30c3",
   32200 => x"0c30c3",
   32201 => x"0c30c3",
   32202 => x"0c30c3",
   32203 => x"0c30c3",
   32204 => x"0c30c3",
   32205 => x"0c30c3",
   32206 => x"0c30c3",
   32207 => x"0c30c3",
   32208 => x"0c30c3",
   32209 => x"0c30c3",
   32210 => x"0c30c3",
   32211 => x"0c30c3",
   32212 => x"0c30c3",
   32213 => x"0c30c3",
   32214 => x"0c30c3",
   32215 => x"0c30c3",
   32216 => x"0c30c3",
   32217 => x"0ebfff",
   32218 => x"ffffff",
   32219 => x"ffffff",
   32220 => x"ffffff",
   32221 => x"ffffff",
   32222 => x"ffffff",
   32223 => x"ffffff",
   32224 => x"ffffff",
   32225 => x"ffffff",
   32226 => x"ffffff",
   32227 => x"ffffff",
   32228 => x"ffffff",
   32229 => x"fffa95",
   32230 => x"abffff",
   32231 => x"ffffff",
   32232 => x"ffffff",
   32233 => x"ffffff",
   32234 => x"ffffff",
   32235 => x"ffffff",
   32236 => x"ffffff",
   32237 => x"ffffff",
   32238 => x"ffffff",
   32239 => x"ffffff",
   32240 => x"ffffff",
   32241 => x"ffffff",
   32242 => x"ffffff",
   32243 => x"ffffff",
   32244 => x"ffffff",
   32245 => x"ffffff",
   32246 => x"ffffff",
   32247 => x"ffffff",
   32248 => x"ffffff",
   32249 => x"ffffff",
   32250 => x"ffffff",
   32251 => x"ffffff",
   32252 => x"ffffff",
   32253 => x"ffffff",
   32254 => x"ffffff",
   32255 => x"ffffff",
   32256 => x"ffffff",
   32257 => x"ffffff",
   32258 => x"ffffff",
   32259 => x"ffffff",
   32260 => x"ffffff",
   32261 => x"ffffff",
   32262 => x"ffffff",
   32263 => x"ffffff",
   32264 => x"ffffff",
   32265 => x"ffffff",
   32266 => x"ffffff",
   32267 => x"ffffff",
   32268 => x"ffffff",
   32269 => x"ffffff",
   32270 => x"ffffff",
   32271 => x"ffffff",
   32272 => x"ffffff",
   32273 => x"ffffff",
   32274 => x"ffffff",
   32275 => x"ffffff",
   32276 => x"ffffff",
   32277 => x"ffffff",
   32278 => x"ffffff",
   32279 => x"ffffff",
   32280 => x"ffffff",
   32281 => x"ffffff",
   32282 => x"ffffff",
   32283 => x"ffffff",
   32284 => x"ffffff",
   32285 => x"ffffff",
   32286 => x"ffffff",
   32287 => x"ffffff",
   32288 => x"ffffff",
   32289 => x"ffffff",
   32290 => x"ffffff",
   32291 => x"ffffff",
   32292 => x"ffffff",
   32293 => x"ffffff",
   32294 => x"ffffff",
   32295 => x"ffffff",
   32296 => x"ffffff",
   32297 => x"ffffff",
   32298 => x"ffffff",
   32299 => x"ffffff",
   32300 => x"ffffff",
   32301 => x"ffffff",
   32302 => x"ffffff",
   32303 => x"ffffff",
   32304 => x"ffffff",
   32305 => x"ffffff",
   32306 => x"ffffff",
   32307 => x"ffffff",
   32308 => x"ffffff",
   32309 => x"ffffff",
   32310 => x"ffffff",
   32311 => x"ffffff",
   32312 => x"ffffff",
   32313 => x"ffffff",
   32314 => x"ffffff",
   32315 => x"ffffff",
   32316 => x"ffffff",
   32317 => x"ffffff",
   32318 => x"ffffff",
   32319 => x"ffffff",
   32320 => x"ffffff",
   32321 => x"ffffff",
   32322 => x"ffffff",
   32323 => x"ffffff",
   32324 => x"ffffff",
   32325 => x"ffffff",
   32326 => x"ffffff",
   32327 => x"ffffff",
   32328 => x"ffffff",
   32329 => x"ffffff",
   32330 => x"ffffff",
   32331 => x"feb0c3",
   32332 => x"0c30c3",
   32333 => x"0c30c3",
   32334 => x"0c30c3",
   32335 => x"0c30c3",
   32336 => x"0c30c3",
   32337 => x"0c30c3",
   32338 => x"0c30c3",
   32339 => x"0c30c3",
   32340 => x"0c30c3",
   32341 => x"0c30c3",
   32342 => x"0c30c3",
   32343 => x"0c30c3",
   32344 => x"0c30c3",
   32345 => x"0c30c3",
   32346 => x"0c30c3",
   32347 => x"0c30c3",
   32348 => x"0c30c3",
   32349 => x"0c30c3",
   32350 => x"0c30c3",
   32351 => x"0c30c3",
   32352 => x"0c30c3",
   32353 => x"0c30c3",
   32354 => x"0c30c3",
   32355 => x"0c30c3",
   32356 => x"0c30c3",
   32357 => x"0c30c3",
   32358 => x"0c30c3",
   32359 => x"0c30c3",
   32360 => x"0c30c3",
   32361 => x"0c30c3",
   32362 => x"0c30c3",
   32363 => x"0c30c3",
   32364 => x"0c30c3",
   32365 => x"0c30c3",
   32366 => x"0c30c3",
   32367 => x"0c30c3",
   32368 => x"0c30c3",
   32369 => x"0c30c3",
   32370 => x"0c30c3",
   32371 => x"0c30c3",
   32372 => x"0c30c3",
   32373 => x"0c30c3",
   32374 => x"0c30c3",
   32375 => x"0c30c3",
   32376 => x"0c30c3",
   32377 => x"5ebfff",
   32378 => x"ffffff",
   32379 => x"ffffff",
   32380 => x"ffffff",
   32381 => x"ffffff",
   32382 => x"ffffff",
   32383 => x"ffffff",
   32384 => x"ffffff",
   32385 => x"ffffff",
   32386 => x"ffffff",
   32387 => x"ffffff",
   32388 => x"ffffff",
   32389 => x"fffa95",
   32390 => x"abffff",
   32391 => x"ffffff",
   32392 => x"ffffff",
   32393 => x"ffffff",
   32394 => x"ffffff",
   32395 => x"ffffff",
   32396 => x"ffffff",
   32397 => x"ffffff",
   32398 => x"ffffff",
   32399 => x"ffffff",
   32400 => x"ffffff",
   32401 => x"ffffff",
   32402 => x"ffffff",
   32403 => x"ffffff",
   32404 => x"ffffff",
   32405 => x"ffffff",
   32406 => x"ffffff",
   32407 => x"ffffff",
   32408 => x"ffffff",
   32409 => x"ffffff",
   32410 => x"ffffff",
   32411 => x"ffffff",
   32412 => x"ffffff",
   32413 => x"ffffff",
   32414 => x"ffffff",
   32415 => x"ffffff",
   32416 => x"ffffff",
   32417 => x"ffffff",
   32418 => x"ffffff",
   32419 => x"ffffff",
   32420 => x"ffffff",
   32421 => x"ffffff",
   32422 => x"ffffff",
   32423 => x"ffffff",
   32424 => x"ffffff",
   32425 => x"ffffff",
   32426 => x"ffffff",
   32427 => x"ffffff",
   32428 => x"ffffff",
   32429 => x"ffffff",
   32430 => x"ffffff",
   32431 => x"ffffff",
   32432 => x"ffffff",
   32433 => x"ffffff",
   32434 => x"ffffff",
   32435 => x"ffffff",
   32436 => x"ffffff",
   32437 => x"ffffff",
   32438 => x"ffffff",
   32439 => x"ffffff",
   32440 => x"ffffff",
   32441 => x"ffffff",
   32442 => x"ffffff",
   32443 => x"ffffff",
   32444 => x"ffffff",
   32445 => x"ffffff",
   32446 => x"ffffff",
   32447 => x"ffffff",
   32448 => x"ffffff",
   32449 => x"ffffff",
   32450 => x"ffffff",
   32451 => x"ffffff",
   32452 => x"ffffff",
   32453 => x"ffffff",
   32454 => x"ffffff",
   32455 => x"ffffff",
   32456 => x"ffffff",
   32457 => x"ffffff",
   32458 => x"ffffff",
   32459 => x"ffffff",
   32460 => x"ffffff",
   32461 => x"ffffff",
   32462 => x"ffffff",
   32463 => x"ffffff",
   32464 => x"ffffff",
   32465 => x"ffffff",
   32466 => x"ffffff",
   32467 => x"ffffff",
   32468 => x"ffffff",
   32469 => x"ffffff",
   32470 => x"ffffff",
   32471 => x"ffffff",
   32472 => x"ffffff",
   32473 => x"ffffff",
   32474 => x"ffffff",
   32475 => x"ffffff",
   32476 => x"ffffff",
   32477 => x"ffffff",
   32478 => x"ffffff",
   32479 => x"ffffff",
   32480 => x"ffffff",
   32481 => x"ffffff",
   32482 => x"ffffff",
   32483 => x"ffffff",
   32484 => x"ffffff",
   32485 => x"ffffff",
   32486 => x"ffffff",
   32487 => x"ffffff",
   32488 => x"ffffff",
   32489 => x"ffffff",
   32490 => x"ffffff",
   32491 => x"feb0c3",
   32492 => x"0c30c3",
   32493 => x"0c30c3",
   32494 => x"0c30c3",
   32495 => x"0c30c3",
   32496 => x"0c30c3",
   32497 => x"0c30c3",
   32498 => x"0c30c3",
   32499 => x"0c30c3",
   32500 => x"0c30c3",
   32501 => x"0c30c3",
   32502 => x"0c30c3",
   32503 => x"0c30c3",
   32504 => x"0c30c3",
   32505 => x"0c30c3",
   32506 => x"0c30c3",
   32507 => x"0c30c3",
   32508 => x"0c30c3",
   32509 => x"0c30c3",
   32510 => x"0c30c3",
   32511 => x"0c30c3",
   32512 => x"0c30c3",
   32513 => x"0c30c3",
   32514 => x"0c30c3",
   32515 => x"0c30c3",
   32516 => x"0c30c3",
   32517 => x"0c30c3",
   32518 => x"0c30c3",
   32519 => x"0c30c3",
   32520 => x"0c30c3",
   32521 => x"0c30c3",
   32522 => x"0c30c3",
   32523 => x"0c30c3",
   32524 => x"0c30c3",
   32525 => x"0c30c3",
   32526 => x"0c30c3",
   32527 => x"0c30c3",
   32528 => x"0c30c3",
   32529 => x"0c30c3",
   32530 => x"0c30c3",
   32531 => x"0c30c3",
   32532 => x"0c30c3",
   32533 => x"0c30c3",
   32534 => x"0c30c3",
   32535 => x"0c30c3",
   32536 => x"0c30c3",
   32537 => x"5ebfff",
   32538 => x"ffffff",
   32539 => x"ffffff",
   32540 => x"ffffff",
   32541 => x"ffffff",
   32542 => x"ffffff",
   32543 => x"ffffff",
   32544 => x"ffffff",
   32545 => x"ffffff",
   32546 => x"ffffff",
   32547 => x"ffffff",
   32548 => x"ffffff",
   32549 => x"fffa95",
   32550 => x"abffff",
   32551 => x"ffffff",
   32552 => x"ffffff",
   32553 => x"ffffff",
   32554 => x"ffffff",
   32555 => x"ffffff",
   32556 => x"ffffff",
   32557 => x"ffffff",
   32558 => x"ffffff",
   32559 => x"ffffff",
   32560 => x"ffffff",
   32561 => x"ffffff",
   32562 => x"ffffff",
   32563 => x"ffffff",
   32564 => x"ffffff",
   32565 => x"ffffff",
   32566 => x"ffffff",
   32567 => x"ffffff",
   32568 => x"ffffff",
   32569 => x"ffffff",
   32570 => x"ffffff",
   32571 => x"ffffff",
   32572 => x"ffffff",
   32573 => x"ffffff",
   32574 => x"ffffff",
   32575 => x"ffffff",
   32576 => x"ffffff",
   32577 => x"ffffff",
   32578 => x"ffffff",
   32579 => x"ffffff",
   32580 => x"ffffff",
   32581 => x"ffffff",
   32582 => x"ffffff",
   32583 => x"ffffff",
   32584 => x"ffffff",
   32585 => x"ffffff",
   32586 => x"ffffff",
   32587 => x"ffffff",
   32588 => x"ffffff",
   32589 => x"ffffff",
   32590 => x"ffffff",
   32591 => x"ffffff",
   32592 => x"ffffff",
   32593 => x"ffffff",
   32594 => x"ffffff",
   32595 => x"ffffff",
   32596 => x"ffffff",
   32597 => x"ffffff",
   32598 => x"ffffff",
   32599 => x"ffffff",
   32600 => x"ffffff",
   32601 => x"ffffff",
   32602 => x"ffffff",
   32603 => x"ffffff",
   32604 => x"ffffff",
   32605 => x"ffffff",
   32606 => x"ffffff",
   32607 => x"ffffff",
   32608 => x"ffffff",
   32609 => x"ffffff",
   32610 => x"ffffff",
   32611 => x"ffffff",
   32612 => x"ffffff",
   32613 => x"ffffff",
   32614 => x"ffffff",
   32615 => x"ffffff",
   32616 => x"ffffff",
   32617 => x"ffffff",
   32618 => x"ffffff",
   32619 => x"ffffff",
   32620 => x"ffffff",
   32621 => x"ffffff",
   32622 => x"ffffff",
   32623 => x"ffffff",
   32624 => x"ffffff",
   32625 => x"ffffff",
   32626 => x"ffffff",
   32627 => x"ffffff",
   32628 => x"ffffff",
   32629 => x"ffffff",
   32630 => x"ffffff",
   32631 => x"ffffff",
   32632 => x"ffffff",
   32633 => x"ffffff",
   32634 => x"ffffff",
   32635 => x"ffffff",
   32636 => x"ffffff",
   32637 => x"ffffff",
   32638 => x"ffffff",
   32639 => x"ffffff",
   32640 => x"ffffff",
   32641 => x"ffffff",
   32642 => x"ffffff",
   32643 => x"ffffff",
   32644 => x"ffffff",
   32645 => x"ffffff",
   32646 => x"ffffff",
   32647 => x"ffffff",
   32648 => x"ffffff",
   32649 => x"ffffff",
   32650 => x"ffffff",
   32651 => x"feb0c3",
   32652 => x"0c30c3",
   32653 => x"0c30c3",
   32654 => x"0c30c3",
   32655 => x"0c30c3",
   32656 => x"0c30c3",
   32657 => x"0c30c3",
   32658 => x"0c30c3",
   32659 => x"0c30c3",
   32660 => x"0c30c3",
   32661 => x"0c30c3",
   32662 => x"0c30c3",
   32663 => x"0c30c3",
   32664 => x"0c30c3",
   32665 => x"0c30c3",
   32666 => x"0c30c3",
   32667 => x"0c30c3",
   32668 => x"0c30c3",
   32669 => x"0c30c3",
   32670 => x"0c30c3",
   32671 => x"0c30c3",
   32672 => x"0c30c3",
   32673 => x"0c30c3",
   32674 => x"0c30c3",
   32675 => x"0c30c3",
   32676 => x"0c30c3",
   32677 => x"0c30c3",
   32678 => x"0c30c3",
   32679 => x"0c30c3",
   32680 => x"0c30c3",
   32681 => x"0c30c3",
   32682 => x"0c30c3",
   32683 => x"0c30c3",
   32684 => x"0c30c3",
   32685 => x"0c30c3",
   32686 => x"0c30c3",
   32687 => x"0c30c3",
   32688 => x"0c30c3",
   32689 => x"0c30c3",
   32690 => x"0c30c3",
   32691 => x"0c30c3",
   32692 => x"0c30c3",
   32693 => x"0c30c3",
   32694 => x"0c30c3",
   32695 => x"0c30c3",
   32696 => x"0c30c3",
   32697 => x"5fffff",
   32698 => x"ffffff",
   32699 => x"ffffff",
   32700 => x"ffffff",
   32701 => x"ffffff",
   32702 => x"ffffff",
   32703 => x"ffffff",
   32704 => x"ffffff",
   32705 => x"ffffff",
   32706 => x"ffffff",
   32707 => x"ffffff",
   32708 => x"ffffff",
   32709 => x"fffa95",
   32710 => x"abffff",
   32711 => x"ffffff",
   32712 => x"ffffff",
   32713 => x"ffffff",
   32714 => x"ffffff",
   32715 => x"ffffff",
   32716 => x"ffffff",
   32717 => x"ffffff",
   32718 => x"ffffff",
   32719 => x"ffffff",
   32720 => x"ffffff",
   32721 => x"ffffff",
   32722 => x"ffffff",
   32723 => x"ffffff",
   32724 => x"ffffff",
   32725 => x"ffffff",
   32726 => x"ffffff",
   32727 => x"ffffff",
   32728 => x"ffffff",
   32729 => x"ffffff",
   32730 => x"ffffff",
   32731 => x"ffffff",
   32732 => x"ffffff",
   32733 => x"ffffff",
   32734 => x"ffffff",
   32735 => x"ffffff",
   32736 => x"ffffff",
   32737 => x"ffffff",
   32738 => x"ffffff",
   32739 => x"ffffff",
   32740 => x"ffffff",
   32741 => x"ffffff",
   32742 => x"ffffff",
   32743 => x"ffffff",
   32744 => x"ffffff",
   32745 => x"ffffff",
   32746 => x"ffffff",
   32747 => x"ffffff",
   32748 => x"ffffff",
   32749 => x"ffffff",
   32750 => x"ffffff",
   32751 => x"ffffff",
   32752 => x"ffffff",
   32753 => x"ffffff",
   32754 => x"ffffff",
   32755 => x"ffffff",
   32756 => x"ffffff",
   32757 => x"ffffff",
   32758 => x"ffffff",
   32759 => x"ffffff",
   32760 => x"ffffff",
   32761 => x"ffffff",
   32762 => x"ffffff",
   32763 => x"ffffff",
   32764 => x"ffffff",
   32765 => x"ffffff",
   32766 => x"ffffff",
   32767 => x"ffffff",
   32768 => x"ffffff",
   32769 => x"ffffff",
   32770 => x"ffffff",
   32771 => x"ffffff",
   32772 => x"ffffff",
   32773 => x"ffffff",
   32774 => x"ffffff",
   32775 => x"ffffff",
   32776 => x"ffffff",
   32777 => x"ffffff",
   32778 => x"ffffff",
   32779 => x"ffffff",
   32780 => x"ffffff",
   32781 => x"ffffff",
   32782 => x"ffffff",
   32783 => x"ffffff",
   32784 => x"ffffff",
   32785 => x"ffffff",
   32786 => x"ffffff",
   32787 => x"ffffff",
   32788 => x"ffffff",
   32789 => x"ffffff",
   32790 => x"ffffff",
   32791 => x"ffffff",
   32792 => x"ffffff",
   32793 => x"ffffff",
   32794 => x"ffffff",
   32795 => x"ffffff",
   32796 => x"ffffff",
   32797 => x"ffffff",
   32798 => x"ffffff",
   32799 => x"ffffff",
   32800 => x"ffffff",
   32801 => x"ffffff",
   32802 => x"ffffff",
   32803 => x"ffffff",
   32804 => x"ffffff",
   32805 => x"ffffff",
   32806 => x"ffffff",
   32807 => x"ffffff",
   32808 => x"ffffff",
   32809 => x"ffffff",
   32810 => x"ffffff",
   32811 => x"feb5c3",
   32812 => x"0c30c3",
   32813 => x"0c30c3",
   32814 => x"0c30c3",
   32815 => x"0c30c3",
   32816 => x"0c30c3",
   32817 => x"0c30c3",
   32818 => x"0c30c3",
   32819 => x"0c30c3",
   32820 => x"0c30c3",
   32821 => x"0c30c3",
   32822 => x"0c30c3",
   32823 => x"0c30c3",
   32824 => x"0c30c3",
   32825 => x"0c30c3",
   32826 => x"0c30c3",
   32827 => x"0c30c3",
   32828 => x"0c30c3",
   32829 => x"0c30c3",
   32830 => x"0c30c3",
   32831 => x"0c30c3",
   32832 => x"0c30c3",
   32833 => x"0c30c3",
   32834 => x"0c30c3",
   32835 => x"0c30c3",
   32836 => x"0c30c3",
   32837 => x"0c30c3",
   32838 => x"0c30c3",
   32839 => x"0c30c3",
   32840 => x"0c30c3",
   32841 => x"0c30c3",
   32842 => x"0c30c3",
   32843 => x"0c30c3",
   32844 => x"0c30c3",
   32845 => x"0c30c3",
   32846 => x"0c30c3",
   32847 => x"0c30c3",
   32848 => x"0c30c3",
   32849 => x"0c30c3",
   32850 => x"0c30c3",
   32851 => x"0c30c3",
   32852 => x"0c30c3",
   32853 => x"0c30c3",
   32854 => x"0c30c3",
   32855 => x"0c30c3",
   32856 => x"0c30c3",
   32857 => x"5fffff",
   32858 => x"ffffff",
   32859 => x"ffffff",
   32860 => x"ffffff",
   32861 => x"ffffff",
   32862 => x"ffffff",
   32863 => x"ffffff",
   32864 => x"ffffff",
   32865 => x"ffffff",
   32866 => x"ffffff",
   32867 => x"ffffff",
   32868 => x"ffffff",
   32869 => x"fffa95",
   32870 => x"abffff",
   32871 => x"ffffff",
   32872 => x"ffffff",
   32873 => x"ffffff",
   32874 => x"ffffff",
   32875 => x"ffffff",
   32876 => x"ffffff",
   32877 => x"ffffff",
   32878 => x"ffffff",
   32879 => x"ffffff",
   32880 => x"ffffff",
   32881 => x"ffffff",
   32882 => x"ffffff",
   32883 => x"ffffff",
   32884 => x"ffffff",
   32885 => x"ffffff",
   32886 => x"ffffff",
   32887 => x"ffffff",
   32888 => x"ffffff",
   32889 => x"ffffff",
   32890 => x"ffffff",
   32891 => x"ffffff",
   32892 => x"ffffff",
   32893 => x"ffffff",
   32894 => x"ffffff",
   32895 => x"ffffff",
   32896 => x"ffffff",
   32897 => x"ffffff",
   32898 => x"ffffff",
   32899 => x"ffffff",
   32900 => x"ffffff",
   32901 => x"ffffff",
   32902 => x"ffffff",
   32903 => x"ffffff",
   32904 => x"ffffff",
   32905 => x"ffffff",
   32906 => x"ffffff",
   32907 => x"ffffff",
   32908 => x"ffffff",
   32909 => x"ffffff",
   32910 => x"ffffff",
   32911 => x"ffffff",
   32912 => x"ffffff",
   32913 => x"ffffff",
   32914 => x"ffffff",
   32915 => x"ffffff",
   32916 => x"ffffff",
   32917 => x"ffffff",
   32918 => x"ffffff",
   32919 => x"ffffff",
   32920 => x"ffffff",
   32921 => x"ffffff",
   32922 => x"ffffff",
   32923 => x"ffffff",
   32924 => x"ffffff",
   32925 => x"ffffff",
   32926 => x"ffffff",
   32927 => x"ffffff",
   32928 => x"ffffff",
   32929 => x"ffffff",
   32930 => x"ffffff",
   32931 => x"ffffff",
   32932 => x"ffffff",
   32933 => x"ffffff",
   32934 => x"ffffff",
   32935 => x"ffffff",
   32936 => x"ffffff",
   32937 => x"ffffff",
   32938 => x"ffffff",
   32939 => x"ffffff",
   32940 => x"ffffff",
   32941 => x"ffffff",
   32942 => x"ffffff",
   32943 => x"ffffff",
   32944 => x"ffffff",
   32945 => x"ffffff",
   32946 => x"ffffff",
   32947 => x"ffffff",
   32948 => x"ffffff",
   32949 => x"ffffff",
   32950 => x"ffffff",
   32951 => x"ffffff",
   32952 => x"ffffff",
   32953 => x"ffffff",
   32954 => x"ffffff",
   32955 => x"ffffff",
   32956 => x"ffffff",
   32957 => x"ffffff",
   32958 => x"ffffff",
   32959 => x"ffffff",
   32960 => x"ffffff",
   32961 => x"ffffff",
   32962 => x"ffffff",
   32963 => x"ffffff",
   32964 => x"ffffff",
   32965 => x"ffffff",
   32966 => x"ffffff",
   32967 => x"ffffff",
   32968 => x"ffffff",
   32969 => x"ffffff",
   32970 => x"ffffff",
   32971 => x"fff5c3",
   32972 => x"0c30c3",
   32973 => x"0c30c3",
   32974 => x"0c30c3",
   32975 => x"0c30c3",
   32976 => x"0c30c3",
   32977 => x"0c30c3",
   32978 => x"0c30c3",
   32979 => x"0c30c3",
   32980 => x"0c30c3",
   32981 => x"0c30c3",
   32982 => x"0c30c3",
   32983 => x"0c30c3",
   32984 => x"0c30c3",
   32985 => x"0c30c3",
   32986 => x"0c30c3",
   32987 => x"0c30c3",
   32988 => x"0c30c3",
   32989 => x"0c30c3",
   32990 => x"0c30c3",
   32991 => x"0c30c3",
   32992 => x"0c30c3",
   32993 => x"0c30c3",
   32994 => x"0c30c3",
   32995 => x"0c30c3",
   32996 => x"0c30c3",
   32997 => x"0c30c3",
   32998 => x"0c30c3",
   32999 => x"0c30c3",
   33000 => x"0c30c3",
   33001 => x"0c30c3",
   33002 => x"0c30c3",
   33003 => x"0c30c3",
   33004 => x"0c30c3",
   33005 => x"0c30c3",
   33006 => x"0c30c3",
   33007 => x"0c30c3",
   33008 => x"0c30c3",
   33009 => x"0c30c3",
   33010 => x"0c30c3",
   33011 => x"0c30c3",
   33012 => x"0c30c3",
   33013 => x"0c30c3",
   33014 => x"0c30c3",
   33015 => x"0c30c3",
   33016 => x"0c30c3",
   33017 => x"5fffff",
   33018 => x"ffffff",
   33019 => x"ffffff",
   33020 => x"ffffff",
   33021 => x"ffffff",
   33022 => x"ffffff",
   33023 => x"ffffff",
   33024 => x"ffffff",
   33025 => x"ffffff",
   33026 => x"ffffff",
   33027 => x"ffffff",
   33028 => x"ffffff",
   33029 => x"fffa95",
   33030 => x"abffff",
   33031 => x"ffffff",
   33032 => x"ffffff",
   33033 => x"ffffff",
   33034 => x"ffffff",
   33035 => x"ffffff",
   33036 => x"ffffff",
   33037 => x"ffffff",
   33038 => x"ffffff",
   33039 => x"ffffff",
   33040 => x"ffffff",
   33041 => x"ffffff",
   33042 => x"ffffff",
   33043 => x"ffffff",
   33044 => x"ffffff",
   33045 => x"ffffff",
   33046 => x"ffffff",
   33047 => x"ffffff",
   33048 => x"ffffff",
   33049 => x"ffffff",
   33050 => x"ffffff",
   33051 => x"ffffff",
   33052 => x"ffffff",
   33053 => x"ffffff",
   33054 => x"ffffff",
   33055 => x"ffffff",
   33056 => x"ffffff",
   33057 => x"ffffff",
   33058 => x"ffffff",
   33059 => x"ffffff",
   33060 => x"ffffff",
   33061 => x"ffffff",
   33062 => x"ffffff",
   33063 => x"ffffff",
   33064 => x"ffffff",
   33065 => x"ffffff",
   33066 => x"ffffff",
   33067 => x"ffffff",
   33068 => x"ffffff",
   33069 => x"ffffff",
   33070 => x"ffffff",
   33071 => x"ffffff",
   33072 => x"ffffff",
   33073 => x"ffffff",
   33074 => x"ffffff",
   33075 => x"ffffff",
   33076 => x"ffffff",
   33077 => x"ffffff",
   33078 => x"ffffff",
   33079 => x"ffffff",
   33080 => x"ffffff",
   33081 => x"ffffff",
   33082 => x"ffffff",
   33083 => x"ffffff",
   33084 => x"ffffff",
   33085 => x"ffffff",
   33086 => x"ffffff",
   33087 => x"ffffff",
   33088 => x"ffffff",
   33089 => x"ffffff",
   33090 => x"ffffff",
   33091 => x"ffffff",
   33092 => x"ffffff",
   33093 => x"ffffff",
   33094 => x"ffffff",
   33095 => x"ffffff",
   33096 => x"ffffff",
   33097 => x"ffffff",
   33098 => x"ffffff",
   33099 => x"ffffff",
   33100 => x"ffffff",
   33101 => x"ffffff",
   33102 => x"ffffff",
   33103 => x"ffffff",
   33104 => x"ffffff",
   33105 => x"ffffff",
   33106 => x"ffffff",
   33107 => x"ffffff",
   33108 => x"ffffff",
   33109 => x"ffffff",
   33110 => x"ffffff",
   33111 => x"ffffff",
   33112 => x"ffffff",
   33113 => x"ffffff",
   33114 => x"ffffff",
   33115 => x"ffffff",
   33116 => x"ffffff",
   33117 => x"ffffff",
   33118 => x"ffffff",
   33119 => x"ffffff",
   33120 => x"ffffff",
   33121 => x"ffffff",
   33122 => x"ffffff",
   33123 => x"ffffff",
   33124 => x"ffffff",
   33125 => x"ffffff",
   33126 => x"ffffff",
   33127 => x"ffffff",
   33128 => x"ffffff",
   33129 => x"ffffff",
   33130 => x"ffffff",
   33131 => x"fff5c3",
   33132 => x"0c30c3",
   33133 => x"0c30c3",
   33134 => x"0c30c3",
   33135 => x"0c30c3",
   33136 => x"0c30c3",
   33137 => x"0c30c3",
   33138 => x"0c30c3",
   33139 => x"0c30c3",
   33140 => x"0c30c3",
   33141 => x"0c30c3",
   33142 => x"0c30c3",
   33143 => x"0c30c3",
   33144 => x"0c30c3",
   33145 => x"0c30c3",
   33146 => x"0c30c3",
   33147 => x"0c30c3",
   33148 => x"0c30c3",
   33149 => x"0c30c3",
   33150 => x"0c30c3",
   33151 => x"0c30c3",
   33152 => x"0c30c3",
   33153 => x"0c30c3",
   33154 => x"0c30c3",
   33155 => x"0c30c3",
   33156 => x"0c30c3",
   33157 => x"0c30c3",
   33158 => x"0c30c3",
   33159 => x"0c30c3",
   33160 => x"0c30c3",
   33161 => x"0c30c3",
   33162 => x"0c30c3",
   33163 => x"0c30c3",
   33164 => x"0c30c3",
   33165 => x"0c30c3",
   33166 => x"0c30c3",
   33167 => x"0c30c3",
   33168 => x"0c30c3",
   33169 => x"0c30c3",
   33170 => x"0c30c3",
   33171 => x"0c30c3",
   33172 => x"0c30c3",
   33173 => x"0c30c3",
   33174 => x"0c30c3",
   33175 => x"0c30c3",
   33176 => x"0c30c3",
   33177 => x"afffff",
   33178 => x"ffffff",
   33179 => x"ffffff",
   33180 => x"ffffff",
   33181 => x"ffffff",
   33182 => x"ffffff",
   33183 => x"ffffff",
   33184 => x"ffffff",
   33185 => x"ffffff",
   33186 => x"ffffff",
   33187 => x"ffffff",
   33188 => x"ffffff",
   33189 => x"fffa95",
   33190 => x"abffff",
   33191 => x"ffffff",
   33192 => x"ffffff",
   33193 => x"ffffff",
   33194 => x"ffffff",
   33195 => x"ffffff",
   33196 => x"ffffff",
   33197 => x"ffffff",
   33198 => x"ffffff",
   33199 => x"ffffff",
   33200 => x"ffffff",
   33201 => x"ffffff",
   33202 => x"ffffff",
   33203 => x"ffffff",
   33204 => x"ffffff",
   33205 => x"ffffff",
   33206 => x"ffffff",
   33207 => x"ffffff",
   33208 => x"ffffff",
   33209 => x"ffffff",
   33210 => x"ffffff",
   33211 => x"ffffff",
   33212 => x"ffffff",
   33213 => x"ffffff",
   33214 => x"ffffff",
   33215 => x"ffffff",
   33216 => x"ffffff",
   33217 => x"ffffff",
   33218 => x"ffffff",
   33219 => x"ffffff",
   33220 => x"ffffff",
   33221 => x"ffffff",
   33222 => x"ffffff",
   33223 => x"ffffff",
   33224 => x"ffffff",
   33225 => x"ffffff",
   33226 => x"ffffff",
   33227 => x"ffffff",
   33228 => x"ffffff",
   33229 => x"ffffff",
   33230 => x"ffffff",
   33231 => x"ffffff",
   33232 => x"ffffff",
   33233 => x"ffffff",
   33234 => x"ffffff",
   33235 => x"ffffff",
   33236 => x"ffffff",
   33237 => x"ffffff",
   33238 => x"ffffff",
   33239 => x"ffffff",
   33240 => x"ffffff",
   33241 => x"ffffff",
   33242 => x"ffffff",
   33243 => x"ffffff",
   33244 => x"ffffff",
   33245 => x"ffffff",
   33246 => x"ffffff",
   33247 => x"ffffff",
   33248 => x"ffffff",
   33249 => x"ffffff",
   33250 => x"ffffff",
   33251 => x"ffffff",
   33252 => x"ffffff",
   33253 => x"ffffff",
   33254 => x"ffffff",
   33255 => x"ffffff",
   33256 => x"ffffff",
   33257 => x"ffffff",
   33258 => x"ffffff",
   33259 => x"ffffff",
   33260 => x"ffffff",
   33261 => x"ffffff",
   33262 => x"ffffff",
   33263 => x"ffffff",
   33264 => x"ffffff",
   33265 => x"ffffff",
   33266 => x"ffffff",
   33267 => x"ffffff",
   33268 => x"ffffff",
   33269 => x"ffffff",
   33270 => x"ffffff",
   33271 => x"ffffff",
   33272 => x"ffffff",
   33273 => x"ffffff",
   33274 => x"ffffff",
   33275 => x"ffffff",
   33276 => x"ffffff",
   33277 => x"ffffff",
   33278 => x"ffffff",
   33279 => x"ffffff",
   33280 => x"ffffff",
   33281 => x"ffffff",
   33282 => x"ffffff",
   33283 => x"ffffff",
   33284 => x"ffffff",
   33285 => x"ffffff",
   33286 => x"ffffff",
   33287 => x"ffffff",
   33288 => x"ffffff",
   33289 => x"ffffff",
   33290 => x"ffffff",
   33291 => x"fffac3",
   33292 => x"0c30c3",
   33293 => x"0c30c3",
   33294 => x"0c30c3",
   33295 => x"0c30c3",
   33296 => x"0c30c3",
   33297 => x"0c30c3",
   33298 => x"0c30c3",
   33299 => x"0c30c3",
   33300 => x"0c30c3",
   33301 => x"0c30c3",
   33302 => x"0c30c3",
   33303 => x"0c30c3",
   33304 => x"0c30c3",
   33305 => x"0c30c3",
   33306 => x"0c30c3",
   33307 => x"0c30c3",
   33308 => x"0c30c3",
   33309 => x"0c30c3",
   33310 => x"0c30c3",
   33311 => x"0c30c3",
   33312 => x"0c30c3",
   33313 => x"0c30c3",
   33314 => x"0c30c3",
   33315 => x"0c30c3",
   33316 => x"0c30c3",
   33317 => x"0c30c3",
   33318 => x"0c30c3",
   33319 => x"0c30c3",
   33320 => x"0c30c3",
   33321 => x"0c30c3",
   33322 => x"0c30c3",
   33323 => x"0c30c3",
   33324 => x"0c30c3",
   33325 => x"0c30c3",
   33326 => x"0c30c3",
   33327 => x"0c30c3",
   33328 => x"0c30c3",
   33329 => x"0c30c3",
   33330 => x"0c30c3",
   33331 => x"0c30c3",
   33332 => x"0c30c3",
   33333 => x"0c30c3",
   33334 => x"0c30c3",
   33335 => x"0c30c3",
   33336 => x"0c30c3",
   33337 => x"afffff",
   33338 => x"ffffff",
   33339 => x"ffffff",
   33340 => x"ffffff",
   33341 => x"ffffff",
   33342 => x"ffffff",
   33343 => x"ffffff",
   33344 => x"ffffff",
   33345 => x"ffffff",
   33346 => x"ffffff",
   33347 => x"ffffff",
   33348 => x"ffffff",
   33349 => x"fffa95",
   33350 => x"abffff",
   33351 => x"ffffff",
   33352 => x"ffffff",
   33353 => x"ffffff",
   33354 => x"ffffff",
   33355 => x"ffffff",
   33356 => x"ffffff",
   33357 => x"ffffff",
   33358 => x"ffffff",
   33359 => x"ffffff",
   33360 => x"ffffff",
   33361 => x"ffffff",
   33362 => x"ffffff",
   33363 => x"ffffff",
   33364 => x"ffffff",
   33365 => x"ffffff",
   33366 => x"ffffff",
   33367 => x"ffffff",
   33368 => x"ffffff",
   33369 => x"ffffff",
   33370 => x"ffffff",
   33371 => x"ffffff",
   33372 => x"ffffff",
   33373 => x"ffffff",
   33374 => x"ffffff",
   33375 => x"ffffff",
   33376 => x"ffffff",
   33377 => x"ffffff",
   33378 => x"ffffff",
   33379 => x"ffffff",
   33380 => x"ffffff",
   33381 => x"ffffff",
   33382 => x"ffffff",
   33383 => x"ffffff",
   33384 => x"ffffff",
   33385 => x"ffffff",
   33386 => x"ffffff",
   33387 => x"ffffff",
   33388 => x"ffffff",
   33389 => x"ffffff",
   33390 => x"ffffff",
   33391 => x"ffffff",
   33392 => x"ffffff",
   33393 => x"ffffff",
   33394 => x"ffffff",
   33395 => x"ffffff",
   33396 => x"ffffff",
   33397 => x"ffffff",
   33398 => x"ffffff",
   33399 => x"ffffff",
   33400 => x"ffffff",
   33401 => x"ffffff",
   33402 => x"ffffff",
   33403 => x"ffffff",
   33404 => x"ffffff",
   33405 => x"ffffff",
   33406 => x"ffffff",
   33407 => x"ffffff",
   33408 => x"ffffff",
   33409 => x"ffffff",
   33410 => x"ffffff",
   33411 => x"ffffff",
   33412 => x"ffffff",
   33413 => x"ffffff",
   33414 => x"ffffff",
   33415 => x"ffffff",
   33416 => x"ffffff",
   33417 => x"ffffff",
   33418 => x"ffffff",
   33419 => x"ffffff",
   33420 => x"ffffff",
   33421 => x"ffffff",
   33422 => x"ffffff",
   33423 => x"ffffff",
   33424 => x"ffffff",
   33425 => x"ffffff",
   33426 => x"ffffff",
   33427 => x"ffffff",
   33428 => x"ffffff",
   33429 => x"ffffff",
   33430 => x"ffffff",
   33431 => x"ffffff",
   33432 => x"ffffff",
   33433 => x"ffffff",
   33434 => x"ffffff",
   33435 => x"ffffff",
   33436 => x"ffffff",
   33437 => x"ffffff",
   33438 => x"ffffff",
   33439 => x"ffffff",
   33440 => x"ffffff",
   33441 => x"ffffff",
   33442 => x"ffffff",
   33443 => x"ffffff",
   33444 => x"ffffff",
   33445 => x"ffffff",
   33446 => x"ffffff",
   33447 => x"ffffff",
   33448 => x"ffffff",
   33449 => x"ffffff",
   33450 => x"ffffff",
   33451 => x"fffac3",
   33452 => x"0c30c3",
   33453 => x"0c30c3",
   33454 => x"0c30c3",
   33455 => x"0c30c3",
   33456 => x"0c30c3",
   33457 => x"0c30c3",
   33458 => x"0c30c3",
   33459 => x"0c30c3",
   33460 => x"0c30c3",
   33461 => x"0c30c3",
   33462 => x"0c30c3",
   33463 => x"0c30c3",
   33464 => x"0c30c3",
   33465 => x"0c30c3",
   33466 => x"0c30c3",
   33467 => x"0c30c3",
   33468 => x"0c30c3",
   33469 => x"0c30c3",
   33470 => x"0c30c3",
   33471 => x"0c30c3",
   33472 => x"0c30c3",
   33473 => x"0c30c3",
   33474 => x"0c30c3",
   33475 => x"0c30c3",
   33476 => x"0c30c3",
   33477 => x"0c30c3",
   33478 => x"0c30c3",
   33479 => x"0c30c3",
   33480 => x"0c30c3",
   33481 => x"0c30c3",
   33482 => x"0c30c3",
   33483 => x"0c30c3",
   33484 => x"0c30c3",
   33485 => x"0c30c3",
   33486 => x"0c30c3",
   33487 => x"0c30c3",
   33488 => x"0c30c3",
   33489 => x"0c30c3",
   33490 => x"0c30c3",
   33491 => x"0c30c3",
   33492 => x"0c30c3",
   33493 => x"0c30c3",
   33494 => x"0c30c3",
   33495 => x"0c30c3",
   33496 => x"0c30d7",
   33497 => x"afffff",
   33498 => x"ffffff",
   33499 => x"ffffff",
   33500 => x"ffffff",
   33501 => x"ffffff",
   33502 => x"ffffff",
   33503 => x"ffffff",
   33504 => x"ffffff",
   33505 => x"ffffff",
   33506 => x"ffffff",
   33507 => x"ffffff",
   33508 => x"ffffff",
   33509 => x"fffa95",
   33510 => x"abffff",
   33511 => x"ffffff",
   33512 => x"ffffff",
   33513 => x"ffffff",
   33514 => x"ffffff",
   33515 => x"ffffff",
   33516 => x"ffffff",
   33517 => x"ffffff",
   33518 => x"ffffff",
   33519 => x"ffffff",
   33520 => x"ffffff",
   33521 => x"ffffff",
   33522 => x"ffffff",
   33523 => x"ffffff",
   33524 => x"ffffff",
   33525 => x"ffffff",
   33526 => x"ffffff",
   33527 => x"ffffff",
   33528 => x"ffffff",
   33529 => x"ffffff",
   33530 => x"ffffff",
   33531 => x"ffffff",
   33532 => x"ffffff",
   33533 => x"ffffff",
   33534 => x"ffffff",
   33535 => x"ffffff",
   33536 => x"ffffff",
   33537 => x"ffffff",
   33538 => x"ffffff",
   33539 => x"ffffff",
   33540 => x"ffffff",
   33541 => x"ffffff",
   33542 => x"ffffff",
   33543 => x"ffffff",
   33544 => x"ffffff",
   33545 => x"ffffff",
   33546 => x"ffffff",
   33547 => x"ffffff",
   33548 => x"ffffff",
   33549 => x"ffffff",
   33550 => x"ffffff",
   33551 => x"ffffff",
   33552 => x"ffffff",
   33553 => x"ffffff",
   33554 => x"ffffff",
   33555 => x"ffffff",
   33556 => x"ffffff",
   33557 => x"ffffff",
   33558 => x"ffffff",
   33559 => x"ffffff",
   33560 => x"ffffff",
   33561 => x"ffffff",
   33562 => x"ffffff",
   33563 => x"ffffff",
   33564 => x"ffffff",
   33565 => x"ffffff",
   33566 => x"ffffff",
   33567 => x"ffffff",
   33568 => x"ffffff",
   33569 => x"ffffff",
   33570 => x"ffffff",
   33571 => x"ffffff",
   33572 => x"ffffff",
   33573 => x"ffffff",
   33574 => x"ffffff",
   33575 => x"ffffff",
   33576 => x"ffffff",
   33577 => x"ffffff",
   33578 => x"ffffff",
   33579 => x"ffffff",
   33580 => x"ffffff",
   33581 => x"ffffff",
   33582 => x"ffffff",
   33583 => x"ffffff",
   33584 => x"ffffff",
   33585 => x"ffffff",
   33586 => x"ffffff",
   33587 => x"ffffff",
   33588 => x"ffffff",
   33589 => x"ffffff",
   33590 => x"ffffff",
   33591 => x"ffffff",
   33592 => x"ffffff",
   33593 => x"ffffff",
   33594 => x"ffffff",
   33595 => x"ffffff",
   33596 => x"ffffff",
   33597 => x"ffffff",
   33598 => x"ffffff",
   33599 => x"ffffff",
   33600 => x"ffffff",
   33601 => x"ffffff",
   33602 => x"ffffff",
   33603 => x"ffffff",
   33604 => x"ffffff",
   33605 => x"ffffff",
   33606 => x"ffffff",
   33607 => x"ffffff",
   33608 => x"ffffff",
   33609 => x"ffffff",
   33610 => x"ffffff",
   33611 => x"fffac3",
   33612 => x"0c30c3",
   33613 => x"0c30c3",
   33614 => x"0c30c3",
   33615 => x"0c30c3",
   33616 => x"0c30c3",
   33617 => x"0c30c3",
   33618 => x"0c30c3",
   33619 => x"0c30c3",
   33620 => x"0c30c3",
   33621 => x"0c30c3",
   33622 => x"0c30c3",
   33623 => x"0c30c3",
   33624 => x"0c30c3",
   33625 => x"0c30c3",
   33626 => x"0c30c3",
   33627 => x"0c30c3",
   33628 => x"0c30c3",
   33629 => x"0c30c3",
   33630 => x"0c30c3",
   33631 => x"0c30c3",
   33632 => x"0c30c3",
   33633 => x"0c30c3",
   33634 => x"0c30c3",
   33635 => x"0c30c3",
   33636 => x"0c30c3",
   33637 => x"0c30c3",
   33638 => x"0c30c3",
   33639 => x"0c30c3",
   33640 => x"0c30c3",
   33641 => x"0c30c3",
   33642 => x"0c30c3",
   33643 => x"0c30c3",
   33644 => x"0c30c3",
   33645 => x"0c30c3",
   33646 => x"0c30c3",
   33647 => x"0c30c3",
   33648 => x"0c30c3",
   33649 => x"0c30c3",
   33650 => x"0c30c3",
   33651 => x"0c30c3",
   33652 => x"0c30c3",
   33653 => x"0c30c3",
   33654 => x"0c30c3",
   33655 => x"0c30c3",
   33656 => x"0c30d7",
   33657 => x"ffffff",
   33658 => x"ffffff",
   33659 => x"ffffff",
   33660 => x"ffffff",
   33661 => x"ffffff",
   33662 => x"ffffff",
   33663 => x"ffffff",
   33664 => x"ffffff",
   33665 => x"ffffff",
   33666 => x"ffffff",
   33667 => x"ffffff",
   33668 => x"ffffff",
   33669 => x"fffa95",
   33670 => x"abffff",
   33671 => x"ffffff",
   33672 => x"ffffff",
   33673 => x"ffffff",
   33674 => x"ffffff",
   33675 => x"ffffff",
   33676 => x"ffffff",
   33677 => x"ffffff",
   33678 => x"ffffff",
   33679 => x"ffffff",
   33680 => x"ffffff",
   33681 => x"ffffff",
   33682 => x"ffffff",
   33683 => x"ffffff",
   33684 => x"ffffff",
   33685 => x"ffffff",
   33686 => x"ffffff",
   33687 => x"ffffff",
   33688 => x"ffffff",
   33689 => x"ffffff",
   33690 => x"ffffff",
   33691 => x"ffffff",
   33692 => x"ffffff",
   33693 => x"ffffff",
   33694 => x"ffffff",
   33695 => x"ffffff",
   33696 => x"ffffff",
   33697 => x"ffffff",
   33698 => x"ffffff",
   33699 => x"ffffff",
   33700 => x"ffffff",
   33701 => x"ffffff",
   33702 => x"ffffff",
   33703 => x"ffffff",
   33704 => x"ffffff",
   33705 => x"ffffff",
   33706 => x"ffffff",
   33707 => x"ffffff",
   33708 => x"ffffff",
   33709 => x"ffffff",
   33710 => x"ffffff",
   33711 => x"ffffff",
   33712 => x"ffffff",
   33713 => x"ffffff",
   33714 => x"ffffff",
   33715 => x"ffffff",
   33716 => x"ffffff",
   33717 => x"ffffff",
   33718 => x"ffffff",
   33719 => x"ffffff",
   33720 => x"ffffff",
   33721 => x"ffffff",
   33722 => x"ffffff",
   33723 => x"ffffff",
   33724 => x"ffffff",
   33725 => x"ffffff",
   33726 => x"ffffff",
   33727 => x"ffffff",
   33728 => x"ffffff",
   33729 => x"ffffff",
   33730 => x"ffffff",
   33731 => x"ffffff",
   33732 => x"ffffff",
   33733 => x"ffffff",
   33734 => x"ffffff",
   33735 => x"ffffff",
   33736 => x"ffffff",
   33737 => x"ffffff",
   33738 => x"ffffff",
   33739 => x"ffffff",
   33740 => x"ffffff",
   33741 => x"ffffff",
   33742 => x"ffffff",
   33743 => x"ffffff",
   33744 => x"ffffff",
   33745 => x"ffffff",
   33746 => x"ffffff",
   33747 => x"ffffff",
   33748 => x"ffffff",
   33749 => x"ffffff",
   33750 => x"ffffff",
   33751 => x"ffffff",
   33752 => x"ffffff",
   33753 => x"ffffff",
   33754 => x"ffffff",
   33755 => x"ffffff",
   33756 => x"ffffff",
   33757 => x"ffffff",
   33758 => x"ffffff",
   33759 => x"ffffff",
   33760 => x"ffffff",
   33761 => x"ffffff",
   33762 => x"ffffff",
   33763 => x"ffffff",
   33764 => x"ffffff",
   33765 => x"ffffff",
   33766 => x"ffffff",
   33767 => x"ffffff",
   33768 => x"ffffff",
   33769 => x"ffffff",
   33770 => x"ffffff",
   33771 => x"fffad7",
   33772 => x"0c30c3",
   33773 => x"0c30c3",
   33774 => x"0c30c3",
   33775 => x"0c30c3",
   33776 => x"0c30c3",
   33777 => x"0c30c3",
   33778 => x"0c30c3",
   33779 => x"0c30c3",
   33780 => x"0c30c3",
   33781 => x"0c30c3",
   33782 => x"0c30c3",
   33783 => x"0c30c3",
   33784 => x"0c30c3",
   33785 => x"0c30c3",
   33786 => x"0c30c3",
   33787 => x"0c30c3",
   33788 => x"0c30c3",
   33789 => x"0c30c3",
   33790 => x"0c30c3",
   33791 => x"0c30c3",
   33792 => x"0c30c3",
   33793 => x"0c30c3",
   33794 => x"0c30c3",
   33795 => x"0c30c3",
   33796 => x"0c30c3",
   33797 => x"0c30c3",
   33798 => x"0c30c3",
   33799 => x"0c30c3",
   33800 => x"0c30c3",
   33801 => x"0c30c3",
   33802 => x"0c30c3",
   33803 => x"0c30c3",
   33804 => x"0c30c3",
   33805 => x"0c30c3",
   33806 => x"0c30c3",
   33807 => x"0c30c3",
   33808 => x"0c30c3",
   33809 => x"0c30c3",
   33810 => x"0c30c3",
   33811 => x"0c30c3",
   33812 => x"0c30c3",
   33813 => x"0c30c3",
   33814 => x"0c30c3",
   33815 => x"0c30c3",
   33816 => x"0c30d7",
   33817 => x"ffffff",
   33818 => x"ffffff",
   33819 => x"ffffff",
   33820 => x"ffffff",
   33821 => x"ffffff",
   33822 => x"ffffff",
   33823 => x"ffffff",
   33824 => x"ffffff",
   33825 => x"ffffff",
   33826 => x"ffffff",
   33827 => x"ffffff",
   33828 => x"ffffff",
   33829 => x"fffa95",
   33830 => x"abffff",
   33831 => x"ffffff",
   33832 => x"ffffff",
   33833 => x"ffffff",
   33834 => x"ffffff",
   33835 => x"ffffff",
   33836 => x"ffffff",
   33837 => x"ffffff",
   33838 => x"ffffff",
   33839 => x"ffffff",
   33840 => x"ffffff",
   33841 => x"ffffff",
   33842 => x"ffffff",
   33843 => x"ffffff",
   33844 => x"ffffff",
   33845 => x"ffffff",
   33846 => x"ffffff",
   33847 => x"ffffff",
   33848 => x"ffffff",
   33849 => x"ffffff",
   33850 => x"ffffff",
   33851 => x"ffffff",
   33852 => x"ffffff",
   33853 => x"ffffff",
   33854 => x"ffffff",
   33855 => x"ffffff",
   33856 => x"ffffff",
   33857 => x"ffffff",
   33858 => x"ffffff",
   33859 => x"ffffff",
   33860 => x"ffffff",
   33861 => x"ffffff",
   33862 => x"ffffff",
   33863 => x"ffffff",
   33864 => x"ffffff",
   33865 => x"ffffff",
   33866 => x"ffffff",
   33867 => x"ffffff",
   33868 => x"ffffff",
   33869 => x"ffffff",
   33870 => x"ffffff",
   33871 => x"ffffff",
   33872 => x"ffffff",
   33873 => x"ffffff",
   33874 => x"ffffff",
   33875 => x"ffffff",
   33876 => x"ffffff",
   33877 => x"ffffff",
   33878 => x"ffffff",
   33879 => x"ffffff",
   33880 => x"ffffff",
   33881 => x"ffffff",
   33882 => x"ffffff",
   33883 => x"ffffff",
   33884 => x"ffffff",
   33885 => x"ffffff",
   33886 => x"ffffff",
   33887 => x"ffffff",
   33888 => x"ffffff",
   33889 => x"ffffff",
   33890 => x"ffffff",
   33891 => x"ffffff",
   33892 => x"ffffff",
   33893 => x"ffffff",
   33894 => x"ffffff",
   33895 => x"ffffff",
   33896 => x"ffffff",
   33897 => x"ffffff",
   33898 => x"ffffff",
   33899 => x"ffffff",
   33900 => x"ffffff",
   33901 => x"ffffff",
   33902 => x"ffffff",
   33903 => x"ffffff",
   33904 => x"ffffff",
   33905 => x"ffffff",
   33906 => x"ffffff",
   33907 => x"ffffff",
   33908 => x"ffffff",
   33909 => x"ffffff",
   33910 => x"ffffff",
   33911 => x"ffffff",
   33912 => x"ffffff",
   33913 => x"ffffff",
   33914 => x"ffffff",
   33915 => x"ffffff",
   33916 => x"ffffff",
   33917 => x"ffffff",
   33918 => x"ffffff",
   33919 => x"ffffff",
   33920 => x"ffffff",
   33921 => x"ffffff",
   33922 => x"ffffff",
   33923 => x"ffffff",
   33924 => x"ffffff",
   33925 => x"ffffff",
   33926 => x"ffffff",
   33927 => x"ffffff",
   33928 => x"ffffff",
   33929 => x"ffffff",
   33930 => x"ffffff",
   33931 => x"ffffd7",
   33932 => x"0c30c3",
   33933 => x"0c30c3",
   33934 => x"0c30c3",
   33935 => x"0c30c3",
   33936 => x"0c30c3",
   33937 => x"0c30c3",
   33938 => x"0c30c3",
   33939 => x"0c30c3",
   33940 => x"0c30c3",
   33941 => x"0c30c3",
   33942 => x"0c30c3",
   33943 => x"0c30c3",
   33944 => x"0c30c3",
   33945 => x"0c30c3",
   33946 => x"0c30c3",
   33947 => x"0c30c3",
   33948 => x"0c30c3",
   33949 => x"0c30c3",
   33950 => x"0c30c3",
   33951 => x"0c30c3",
   33952 => x"0c30c3",
   33953 => x"0c30c3",
   33954 => x"0c30c3",
   33955 => x"0c30c3",
   33956 => x"0c30c3",
   33957 => x"0c30c3",
   33958 => x"0c30c3",
   33959 => x"0c30c3",
   33960 => x"0c30c3",
   33961 => x"0c30c3",
   33962 => x"0c30c3",
   33963 => x"0c30c3",
   33964 => x"0c30c3",
   33965 => x"0c30c3",
   33966 => x"0c30c3",
   33967 => x"0c30c3",
   33968 => x"0c30c3",
   33969 => x"0c30c3",
   33970 => x"0c30c3",
   33971 => x"0c30c3",
   33972 => x"0c30c3",
   33973 => x"0c30c3",
   33974 => x"0c30c3",
   33975 => x"0c30c3",
   33976 => x"0c30eb",
   33977 => x"ffffff",
   33978 => x"ffffff",
   33979 => x"ffffff",
   33980 => x"ffffff",
   33981 => x"ffffff",
   33982 => x"ffffff",
   33983 => x"ffffff",
   33984 => x"ffffff",
   33985 => x"ffffff",
   33986 => x"ffffff",
   33987 => x"ffffff",
   33988 => x"ffffff",
   33989 => x"fffa95",
   33990 => x"abffff",
   33991 => x"ffffff",
   33992 => x"ffffff",
   33993 => x"ffffff",
   33994 => x"ffffff",
   33995 => x"ffffff",
   33996 => x"ffffff",
   33997 => x"ffffff",
   33998 => x"ffffff",
   33999 => x"ffffff",
   34000 => x"ffffff",
   34001 => x"ffffff",
   34002 => x"ffffff",
   34003 => x"ffffff",
   34004 => x"ffffff",
   34005 => x"ffffff",
   34006 => x"ffffff",
   34007 => x"ffffff",
   34008 => x"ffffff",
   34009 => x"ffffff",
   34010 => x"ffffff",
   34011 => x"ffffff",
   34012 => x"ffffff",
   34013 => x"ffffff",
   34014 => x"ffffff",
   34015 => x"ffffff",
   34016 => x"ffffff",
   34017 => x"ffffff",
   34018 => x"ffffff",
   34019 => x"ffffff",
   34020 => x"ffffff",
   34021 => x"ffffff",
   34022 => x"ffffff",
   34023 => x"ffffff",
   34024 => x"ffffff",
   34025 => x"ffffff",
   34026 => x"ffffff",
   34027 => x"ffffff",
   34028 => x"ffffff",
   34029 => x"ffffff",
   34030 => x"ffffff",
   34031 => x"ffffff",
   34032 => x"ffffff",
   34033 => x"ffffff",
   34034 => x"ffffff",
   34035 => x"ffffff",
   34036 => x"ffffff",
   34037 => x"ffffff",
   34038 => x"ffffff",
   34039 => x"ffffff",
   34040 => x"ffffff",
   34041 => x"ffffff",
   34042 => x"ffffff",
   34043 => x"ffffff",
   34044 => x"ffffff",
   34045 => x"ffffff",
   34046 => x"ffffff",
   34047 => x"ffffff",
   34048 => x"ffffff",
   34049 => x"ffffff",
   34050 => x"ffffff",
   34051 => x"ffffff",
   34052 => x"ffffff",
   34053 => x"ffffff",
   34054 => x"ffffff",
   34055 => x"ffffff",
   34056 => x"ffffff",
   34057 => x"ffffff",
   34058 => x"ffffff",
   34059 => x"ffffff",
   34060 => x"ffffff",
   34061 => x"ffffff",
   34062 => x"ffffff",
   34063 => x"ffffff",
   34064 => x"ffffff",
   34065 => x"ffffff",
   34066 => x"ffffff",
   34067 => x"ffffff",
   34068 => x"ffffff",
   34069 => x"ffffff",
   34070 => x"ffffff",
   34071 => x"ffffff",
   34072 => x"ffffff",
   34073 => x"ffffff",
   34074 => x"ffffff",
   34075 => x"ffffff",
   34076 => x"ffffff",
   34077 => x"ffffff",
   34078 => x"ffffff",
   34079 => x"ffffff",
   34080 => x"ffffff",
   34081 => x"ffffff",
   34082 => x"ffffff",
   34083 => x"ffffff",
   34084 => x"ffffff",
   34085 => x"ffffff",
   34086 => x"ffffff",
   34087 => x"ffffff",
   34088 => x"ffffff",
   34089 => x"ffffff",
   34090 => x"ffffff",
   34091 => x"ffffeb",
   34092 => x"0c30c3",
   34093 => x"0c30c3",
   34094 => x"0c30c3",
   34095 => x"0c30c3",
   34096 => x"0c30c3",
   34097 => x"0c30c3",
   34098 => x"0c30c3",
   34099 => x"0c30c3",
   34100 => x"0c30c3",
   34101 => x"0c30c3",
   34102 => x"0c30c3",
   34103 => x"0c30c3",
   34104 => x"0c30c3",
   34105 => x"0c30c3",
   34106 => x"0c30c3",
   34107 => x"0c30c3",
   34108 => x"0c30c3",
   34109 => x"0c30c3",
   34110 => x"0c30c3",
   34111 => x"0c30c3",
   34112 => x"0c30c3",
   34113 => x"0c30c3",
   34114 => x"0c30c3",
   34115 => x"0c30c3",
   34116 => x"0c30c3",
   34117 => x"0c30c3",
   34118 => x"0c30c3",
   34119 => x"0c30c3",
   34120 => x"0c30c3",
   34121 => x"0c30c3",
   34122 => x"0c30c3",
   34123 => x"0c30c3",
   34124 => x"0c30c3",
   34125 => x"0c30c3",
   34126 => x"0c30c3",
   34127 => x"0c30c3",
   34128 => x"0c30c3",
   34129 => x"0c30c3",
   34130 => x"0c30c3",
   34131 => x"0c30c3",
   34132 => x"0c30c3",
   34133 => x"0c30c3",
   34134 => x"0c30c3",
   34135 => x"0c30c3",
   34136 => x"0c35eb",
   34137 => x"ffffff",
   34138 => x"ffffff",
   34139 => x"ffffff",
   34140 => x"ffffff",
   34141 => x"ffffff",
   34142 => x"ffffff",
   34143 => x"ffffff",
   34144 => x"ffffff",
   34145 => x"ffffff",
   34146 => x"ffffff",
   34147 => x"ffffff",
   34148 => x"ffffff",
   34149 => x"fffa95",
   34150 => x"abffff",
   34151 => x"ffffff",
   34152 => x"ffffff",
   34153 => x"ffffff",
   34154 => x"ffffff",
   34155 => x"ffffff",
   34156 => x"ffffff",
   34157 => x"ffffff",
   34158 => x"ffffff",
   34159 => x"ffffff",
   34160 => x"ffffff",
   34161 => x"ffffff",
   34162 => x"ffffff",
   34163 => x"ffffff",
   34164 => x"ffffff",
   34165 => x"ffffff",
   34166 => x"ffffff",
   34167 => x"ffffff",
   34168 => x"ffffff",
   34169 => x"ffffff",
   34170 => x"ffffff",
   34171 => x"ffffff",
   34172 => x"ffffff",
   34173 => x"ffffff",
   34174 => x"ffffff",
   34175 => x"ffffff",
   34176 => x"ffffff",
   34177 => x"ffffff",
   34178 => x"ffffff",
   34179 => x"ffffff",
   34180 => x"ffffff",
   34181 => x"ffffff",
   34182 => x"ffffff",
   34183 => x"ffffff",
   34184 => x"ffffff",
   34185 => x"ffffff",
   34186 => x"ffffff",
   34187 => x"ffffff",
   34188 => x"ffffff",
   34189 => x"ffffff",
   34190 => x"ffffff",
   34191 => x"ffffff",
   34192 => x"ffffff",
   34193 => x"ffffff",
   34194 => x"ffffff",
   34195 => x"ffffff",
   34196 => x"ffffff",
   34197 => x"ffffff",
   34198 => x"ffffff",
   34199 => x"ffffff",
   34200 => x"ffffff",
   34201 => x"ffffff",
   34202 => x"ffffff",
   34203 => x"ffffff",
   34204 => x"ffffff",
   34205 => x"ffffff",
   34206 => x"ffffff",
   34207 => x"ffffff",
   34208 => x"ffffff",
   34209 => x"ffffff",
   34210 => x"ffffff",
   34211 => x"ffffff",
   34212 => x"ffffff",
   34213 => x"ffffff",
   34214 => x"ffffff",
   34215 => x"ffffff",
   34216 => x"ffffff",
   34217 => x"ffffff",
   34218 => x"ffffff",
   34219 => x"ffffff",
   34220 => x"ffffff",
   34221 => x"ffffff",
   34222 => x"ffffff",
   34223 => x"ffffff",
   34224 => x"ffffff",
   34225 => x"ffffff",
   34226 => x"ffffff",
   34227 => x"ffffff",
   34228 => x"ffffff",
   34229 => x"ffffff",
   34230 => x"ffffff",
   34231 => x"ffffff",
   34232 => x"ffffff",
   34233 => x"ffffff",
   34234 => x"ffffff",
   34235 => x"ffffff",
   34236 => x"ffffff",
   34237 => x"ffffff",
   34238 => x"ffffff",
   34239 => x"ffffff",
   34240 => x"ffffff",
   34241 => x"ffffff",
   34242 => x"ffffff",
   34243 => x"ffffff",
   34244 => x"ffffff",
   34245 => x"ffffff",
   34246 => x"ffffff",
   34247 => x"ffffff",
   34248 => x"ffffff",
   34249 => x"ffffff",
   34250 => x"ffffff",
   34251 => x"ffffeb",
   34252 => x"0c30c3",
   34253 => x"0c30c3",
   34254 => x"0c30c3",
   34255 => x"0c30c3",
   34256 => x"0c30c3",
   34257 => x"0c30c3",
   34258 => x"0c30c3",
   34259 => x"0c30c3",
   34260 => x"0c30c3",
   34261 => x"0c30c3",
   34262 => x"0c30c3",
   34263 => x"0c30c3",
   34264 => x"0c30c3",
   34265 => x"0c30c3",
   34266 => x"0c30c3",
   34267 => x"0c30c3",
   34268 => x"0c30c3",
   34269 => x"0c30c3",
   34270 => x"0c30c3",
   34271 => x"0c30c3",
   34272 => x"0c30c3",
   34273 => x"0c30c3",
   34274 => x"0c30c3",
   34275 => x"0c30c3",
   34276 => x"0c30c3",
   34277 => x"0c30c3",
   34278 => x"0c30c3",
   34279 => x"0c30c3",
   34280 => x"0c30c3",
   34281 => x"0c30c3",
   34282 => x"0c30c3",
   34283 => x"0c30c3",
   34284 => x"0c30c3",
   34285 => x"0c30c3",
   34286 => x"0c30c3",
   34287 => x"0c30c3",
   34288 => x"0c30c3",
   34289 => x"0c30c3",
   34290 => x"0c30c3",
   34291 => x"0c30c3",
   34292 => x"0c30c3",
   34293 => x"0c30c3",
   34294 => x"0c30c3",
   34295 => x"0c30c3",
   34296 => x"0c35ff",
   34297 => x"ffffff",
   34298 => x"ffffff",
   34299 => x"ffffff",
   34300 => x"ffffff",
   34301 => x"ffffff",
   34302 => x"ffffff",
   34303 => x"ffffff",
   34304 => x"ffffff",
   34305 => x"ffffff",
   34306 => x"ffffff",
   34307 => x"ffffff",
   34308 => x"ffffff",
   34309 => x"fffa95",
   34310 => x"abffff",
   34311 => x"ffffff",
   34312 => x"ffffff",
   34313 => x"ffffff",
   34314 => x"ffffff",
   34315 => x"ffffff",
   34316 => x"ffffff",
   34317 => x"ffffff",
   34318 => x"ffffff",
   34319 => x"ffffff",
   34320 => x"ffffff",
   34321 => x"ffffff",
   34322 => x"ffffff",
   34323 => x"ffffff",
   34324 => x"ffffff",
   34325 => x"ffffff",
   34326 => x"ffffff",
   34327 => x"ffffff",
   34328 => x"ffffff",
   34329 => x"ffffff",
   34330 => x"ffffff",
   34331 => x"ffffff",
   34332 => x"ffffff",
   34333 => x"ffffff",
   34334 => x"ffffff",
   34335 => x"ffffff",
   34336 => x"ffffff",
   34337 => x"ffffff",
   34338 => x"ffffff",
   34339 => x"ffffff",
   34340 => x"ffffff",
   34341 => x"ffffff",
   34342 => x"ffffff",
   34343 => x"ffffff",
   34344 => x"ffffff",
   34345 => x"ffffff",
   34346 => x"ffffff",
   34347 => x"ffffff",
   34348 => x"ffffff",
   34349 => x"ffffff",
   34350 => x"ffffff",
   34351 => x"ffffff",
   34352 => x"ffffff",
   34353 => x"ffffff",
   34354 => x"ffffff",
   34355 => x"ffffff",
   34356 => x"ffffff",
   34357 => x"ffffff",
   34358 => x"ffffff",
   34359 => x"ffffff",
   34360 => x"ffffff",
   34361 => x"ffffff",
   34362 => x"ffffff",
   34363 => x"ffffff",
   34364 => x"ffffff",
   34365 => x"ffffff",
   34366 => x"ffffff",
   34367 => x"ffffff",
   34368 => x"ffffff",
   34369 => x"ffffff",
   34370 => x"ffffff",
   34371 => x"ffffff",
   34372 => x"ffffff",
   34373 => x"ffffff",
   34374 => x"ffffff",
   34375 => x"ffffff",
   34376 => x"ffffff",
   34377 => x"ffffff",
   34378 => x"ffffff",
   34379 => x"ffffff",
   34380 => x"ffffff",
   34381 => x"ffffff",
   34382 => x"ffffff",
   34383 => x"ffffff",
   34384 => x"ffffff",
   34385 => x"ffffff",
   34386 => x"ffffff",
   34387 => x"ffffff",
   34388 => x"ffffff",
   34389 => x"ffffff",
   34390 => x"ffffff",
   34391 => x"ffffff",
   34392 => x"ffffff",
   34393 => x"ffffff",
   34394 => x"ffffff",
   34395 => x"ffffff",
   34396 => x"ffffff",
   34397 => x"ffffff",
   34398 => x"ffffff",
   34399 => x"ffffff",
   34400 => x"ffffff",
   34401 => x"ffffff",
   34402 => x"ffffff",
   34403 => x"ffffff",
   34404 => x"ffffff",
   34405 => x"ffffff",
   34406 => x"ffffff",
   34407 => x"ffffff",
   34408 => x"ffffff",
   34409 => x"ffffff",
   34410 => x"ffffff",
   34411 => x"ffffff",
   34412 => x"5c30c3",
   34413 => x"0c30c3",
   34414 => x"0c30c3",
   34415 => x"0c30c3",
   34416 => x"0c30c3",
   34417 => x"0c30c3",
   34418 => x"0c30c3",
   34419 => x"0c30c3",
   34420 => x"0c30c3",
   34421 => x"0c30c3",
   34422 => x"0c30c3",
   34423 => x"0c30c3",
   34424 => x"0c30c3",
   34425 => x"0c30c3",
   34426 => x"0c30c3",
   34427 => x"0c30c3",
   34428 => x"0c30c3",
   34429 => x"0c30c3",
   34430 => x"0c30c3",
   34431 => x"0c30c3",
   34432 => x"0c30c3",
   34433 => x"0c30c3",
   34434 => x"0c30c3",
   34435 => x"0c30c3",
   34436 => x"0c30c3",
   34437 => x"0c30c3",
   34438 => x"0c30c3",
   34439 => x"0c30c3",
   34440 => x"0c30c3",
   34441 => x"0c30c3",
   34442 => x"0c30c3",
   34443 => x"0c30c3",
   34444 => x"0c30c3",
   34445 => x"0c30c3",
   34446 => x"0c30c3",
   34447 => x"0c30c3",
   34448 => x"0c30c3",
   34449 => x"0c30c3",
   34450 => x"0c30c3",
   34451 => x"0c30c3",
   34452 => x"0c30c3",
   34453 => x"0c30c3",
   34454 => x"0c30c3",
   34455 => x"0c30c3",
   34456 => x"0c35ff",
   34457 => x"ffffff",
   34458 => x"ffffff",
   34459 => x"ffffff",
   34460 => x"ffffff",
   34461 => x"ffffff",
   34462 => x"ffffff",
   34463 => x"ffffff",
   34464 => x"ffffff",
   34465 => x"ffffff",
   34466 => x"ffffff",
   34467 => x"ffffff",
   34468 => x"ffffff",
   34469 => x"fffa95",
   34470 => x"abffff",
   34471 => x"ffffff",
   34472 => x"ffffff",
   34473 => x"ffffff",
   34474 => x"ffffff",
   34475 => x"ffffff",
   34476 => x"ffffff",
   34477 => x"ffffff",
   34478 => x"ffffff",
   34479 => x"ffffff",
   34480 => x"ffffff",
   34481 => x"ffffff",
   34482 => x"ffffff",
   34483 => x"ffffff",
   34484 => x"ffffff",
   34485 => x"ffffff",
   34486 => x"ffffff",
   34487 => x"ffffff",
   34488 => x"ffffff",
   34489 => x"ffffff",
   34490 => x"ffffff",
   34491 => x"ffffff",
   34492 => x"ffffff",
   34493 => x"ffffff",
   34494 => x"ffffff",
   34495 => x"ffffff",
   34496 => x"ffffff",
   34497 => x"ffffff",
   34498 => x"ffffff",
   34499 => x"ffffff",
   34500 => x"ffffff",
   34501 => x"ffffff",
   34502 => x"ffffff",
   34503 => x"ffffff",
   34504 => x"ffffff",
   34505 => x"ffffff",
   34506 => x"ffffff",
   34507 => x"ffffff",
   34508 => x"ffffff",
   34509 => x"ffffff",
   34510 => x"ffffff",
   34511 => x"ffffff",
   34512 => x"ffffff",
   34513 => x"ffffff",
   34514 => x"ffffff",
   34515 => x"ffffff",
   34516 => x"ffffff",
   34517 => x"ffffff",
   34518 => x"ffffff",
   34519 => x"ffffff",
   34520 => x"ffffff",
   34521 => x"ffffff",
   34522 => x"ffffff",
   34523 => x"ffffff",
   34524 => x"ffffff",
   34525 => x"ffffff",
   34526 => x"ffffff",
   34527 => x"ffffff",
   34528 => x"ffffff",
   34529 => x"ffffff",
   34530 => x"ffffff",
   34531 => x"ffffff",
   34532 => x"ffffff",
   34533 => x"ffffff",
   34534 => x"ffffff",
   34535 => x"ffffff",
   34536 => x"ffffff",
   34537 => x"ffffff",
   34538 => x"ffffff",
   34539 => x"ffffff",
   34540 => x"ffffff",
   34541 => x"ffffff",
   34542 => x"ffffff",
   34543 => x"ffffff",
   34544 => x"ffffff",
   34545 => x"ffffff",
   34546 => x"ffffff",
   34547 => x"ffffff",
   34548 => x"ffffff",
   34549 => x"ffffff",
   34550 => x"ffffff",
   34551 => x"ffffff",
   34552 => x"ffffff",
   34553 => x"ffffff",
   34554 => x"ffffff",
   34555 => x"ffffff",
   34556 => x"ffffff",
   34557 => x"ffffff",
   34558 => x"ffffff",
   34559 => x"ffffff",
   34560 => x"ffffff",
   34561 => x"ffffff",
   34562 => x"ffffff",
   34563 => x"ffffff",
   34564 => x"ffffff",
   34565 => x"ffffff",
   34566 => x"ffffff",
   34567 => x"ffffff",
   34568 => x"ffffff",
   34569 => x"ffffff",
   34570 => x"ffffff",
   34571 => x"ffffff",
   34572 => x"5c30c3",
   34573 => x"0c30c3",
   34574 => x"0c30c3",
   34575 => x"0c30c3",
   34576 => x"0c30c3",
   34577 => x"0c30c3",
   34578 => x"0c30c3",
   34579 => x"0c30c3",
   34580 => x"0c30c3",
   34581 => x"0c30c3",
   34582 => x"0c30c3",
   34583 => x"0c30c3",
   34584 => x"0c30c3",
   34585 => x"0c30c3",
   34586 => x"0c30c3",
   34587 => x"0c30c3",
   34588 => x"0c30c3",
   34589 => x"0c30c3",
   34590 => x"0c30c3",
   34591 => x"0c30c3",
   34592 => x"0c30c3",
   34593 => x"0c30c3",
   34594 => x"0c30c3",
   34595 => x"0c30c3",
   34596 => x"0c30c3",
   34597 => x"0c30c3",
   34598 => x"0c30c3",
   34599 => x"0c30c3",
   34600 => x"0c30c3",
   34601 => x"0c30c3",
   34602 => x"0c30c3",
   34603 => x"0c30c3",
   34604 => x"0c30c3",
   34605 => x"0c30c3",
   34606 => x"0c30c3",
   34607 => x"0c30c3",
   34608 => x"0c30c3",
   34609 => x"0c30c3",
   34610 => x"0c30c3",
   34611 => x"0c30c3",
   34612 => x"0c30c3",
   34613 => x"0c30c3",
   34614 => x"0c30c3",
   34615 => x"0c30c3",
   34616 => x"0c3aff",
   34617 => x"ffffff",
   34618 => x"ffffff",
   34619 => x"ffffff",
   34620 => x"ffffff",
   34621 => x"ffffff",
   34622 => x"ffffff",
   34623 => x"ffffff",
   34624 => x"ffffff",
   34625 => x"ffffff",
   34626 => x"ffffff",
   34627 => x"ffffff",
   34628 => x"ffffff",
   34629 => x"fffa95",
   34630 => x"abffff",
   34631 => x"ffffff",
   34632 => x"ffffff",
   34633 => x"ffffff",
   34634 => x"ffffff",
   34635 => x"ffffff",
   34636 => x"ffffff",
   34637 => x"ffffff",
   34638 => x"ffffff",
   34639 => x"ffffff",
   34640 => x"ffffff",
   34641 => x"ffffff",
   34642 => x"ffffff",
   34643 => x"ffffff",
   34644 => x"ffffff",
   34645 => x"ffffff",
   34646 => x"ffffff",
   34647 => x"ffffff",
   34648 => x"ffffff",
   34649 => x"ffffff",
   34650 => x"ffffff",
   34651 => x"ffffff",
   34652 => x"ffffff",
   34653 => x"ffffff",
   34654 => x"ffffff",
   34655 => x"ffffff",
   34656 => x"ffffff",
   34657 => x"ffffff",
   34658 => x"ffffff",
   34659 => x"ffffff",
   34660 => x"ffffff",
   34661 => x"ffffff",
   34662 => x"ffffff",
   34663 => x"ffffff",
   34664 => x"ffffff",
   34665 => x"ffffff",
   34666 => x"ffffff",
   34667 => x"ffffff",
   34668 => x"ffffff",
   34669 => x"ffffff",
   34670 => x"ffffff",
   34671 => x"ffffff",
   34672 => x"ffffff",
   34673 => x"ffffff",
   34674 => x"ffffff",
   34675 => x"ffffff",
   34676 => x"ffffff",
   34677 => x"ffffff",
   34678 => x"ffffff",
   34679 => x"ffffff",
   34680 => x"ffffff",
   34681 => x"ffffff",
   34682 => x"ffffff",
   34683 => x"ffffff",
   34684 => x"ffffff",
   34685 => x"ffffff",
   34686 => x"ffffff",
   34687 => x"ffffff",
   34688 => x"ffffff",
   34689 => x"ffffff",
   34690 => x"ffffff",
   34691 => x"ffffff",
   34692 => x"ffffff",
   34693 => x"ffffff",
   34694 => x"ffffff",
   34695 => x"ffffff",
   34696 => x"ffffff",
   34697 => x"ffffff",
   34698 => x"ffffff",
   34699 => x"ffffff",
   34700 => x"ffffff",
   34701 => x"ffffff",
   34702 => x"ffffff",
   34703 => x"ffffff",
   34704 => x"ffffff",
   34705 => x"ffffff",
   34706 => x"ffffff",
   34707 => x"ffffff",
   34708 => x"ffffff",
   34709 => x"ffffff",
   34710 => x"ffffff",
   34711 => x"ffffff",
   34712 => x"ffffff",
   34713 => x"ffffff",
   34714 => x"ffffff",
   34715 => x"ffffff",
   34716 => x"ffffff",
   34717 => x"ffffff",
   34718 => x"ffffff",
   34719 => x"ffffff",
   34720 => x"ffffff",
   34721 => x"ffffff",
   34722 => x"ffffff",
   34723 => x"ffffff",
   34724 => x"ffffff",
   34725 => x"ffffff",
   34726 => x"ffffff",
   34727 => x"ffffff",
   34728 => x"ffffff",
   34729 => x"ffffff",
   34730 => x"ffffff",
   34731 => x"ffffff",
   34732 => x"ac30c3",
   34733 => x"0c30c3",
   34734 => x"0c30c3",
   34735 => x"0c30c3",
   34736 => x"0c30c3",
   34737 => x"0c30c3",
   34738 => x"0c30c3",
   34739 => x"0c30c3",
   34740 => x"0c30c3",
   34741 => x"0c30c3",
   34742 => x"0c30c3",
   34743 => x"0c30c3",
   34744 => x"0c30c3",
   34745 => x"0c30c3",
   34746 => x"0c30c3",
   34747 => x"0c30c3",
   34748 => x"0c30c3",
   34749 => x"0c30c3",
   34750 => x"0c30c3",
   34751 => x"0c30c3",
   34752 => x"0c30c3",
   34753 => x"0c30c3",
   34754 => x"0c30c3",
   34755 => x"0c30c3",
   34756 => x"0c30c3",
   34757 => x"0c30c3",
   34758 => x"0c30c3",
   34759 => x"0c30c3",
   34760 => x"0c30c3",
   34761 => x"0c30c3",
   34762 => x"0c30c3",
   34763 => x"0c30c3",
   34764 => x"0c30c3",
   34765 => x"0c30c3",
   34766 => x"0c30c3",
   34767 => x"0c30c3",
   34768 => x"0c30c3",
   34769 => x"0c30c3",
   34770 => x"0c30c3",
   34771 => x"0c30c3",
   34772 => x"0c30c3",
   34773 => x"0c30c3",
   34774 => x"0c30c3",
   34775 => x"0c30c3",
   34776 => x"0d7aff",
   34777 => x"ffffff",
   34778 => x"ffffff",
   34779 => x"ffffff",
   34780 => x"ffffff",
   34781 => x"ffffff",
   34782 => x"ffffff",
   34783 => x"ffffff",
   34784 => x"ffffff",
   34785 => x"ffffff",
   34786 => x"ffffff",
   34787 => x"ffffff",
   34788 => x"ffffff",
   34789 => x"fffa95",
   34790 => x"abffff",
   34791 => x"ffffff",
   34792 => x"ffffff",
   34793 => x"ffffff",
   34794 => x"ffffff",
   34795 => x"ffffff",
   34796 => x"ffffff",
   34797 => x"ffffff",
   34798 => x"ffffff",
   34799 => x"ffffff",
   34800 => x"ffffff",
   34801 => x"ffffff",
   34802 => x"ffffff",
   34803 => x"ffffff",
   34804 => x"ffffff",
   34805 => x"ffffff",
   34806 => x"ffffff",
   34807 => x"ffffff",
   34808 => x"ffffff",
   34809 => x"ffffff",
   34810 => x"ffffff",
   34811 => x"ffffff",
   34812 => x"ffffff",
   34813 => x"ffffff",
   34814 => x"ffffff",
   34815 => x"ffffff",
   34816 => x"ffffff",
   34817 => x"ffffff",
   34818 => x"ffffff",
   34819 => x"ffffff",
   34820 => x"ffffff",
   34821 => x"ffffff",
   34822 => x"ffffff",
   34823 => x"ffffff",
   34824 => x"ffffff",
   34825 => x"ffffff",
   34826 => x"ffffff",
   34827 => x"ffffff",
   34828 => x"ffffff",
   34829 => x"ffffff",
   34830 => x"ffffff",
   34831 => x"ffffff",
   34832 => x"ffffff",
   34833 => x"ffffff",
   34834 => x"ffffff",
   34835 => x"ffffff",
   34836 => x"ffffff",
   34837 => x"ffffff",
   34838 => x"ffffff",
   34839 => x"ffffff",
   34840 => x"ffffff",
   34841 => x"ffffff",
   34842 => x"ffffff",
   34843 => x"ffffff",
   34844 => x"ffffff",
   34845 => x"ffffff",
   34846 => x"ffffff",
   34847 => x"ffffff",
   34848 => x"ffffff",
   34849 => x"ffffff",
   34850 => x"ffffff",
   34851 => x"ffffff",
   34852 => x"ffffff",
   34853 => x"ffffff",
   34854 => x"ffffff",
   34855 => x"ffffff",
   34856 => x"ffffff",
   34857 => x"ffffff",
   34858 => x"ffffff",
   34859 => x"ffffff",
   34860 => x"ffffff",
   34861 => x"ffffff",
   34862 => x"ffffff",
   34863 => x"ffffff",
   34864 => x"ffffff",
   34865 => x"ffffff",
   34866 => x"ffffff",
   34867 => x"ffffff",
   34868 => x"ffffff",
   34869 => x"ffffff",
   34870 => x"ffffff",
   34871 => x"ffffff",
   34872 => x"ffffff",
   34873 => x"ffffff",
   34874 => x"ffffff",
   34875 => x"ffffff",
   34876 => x"ffffff",
   34877 => x"ffffff",
   34878 => x"ffffff",
   34879 => x"ffffff",
   34880 => x"ffffff",
   34881 => x"ffffff",
   34882 => x"ffffff",
   34883 => x"ffffff",
   34884 => x"ffffff",
   34885 => x"ffffff",
   34886 => x"ffffff",
   34887 => x"ffffff",
   34888 => x"ffffff",
   34889 => x"ffffff",
   34890 => x"ffffff",
   34891 => x"ffffff",
   34892 => x"ac30c3",
   34893 => x"0c30c3",
   34894 => x"0c30c3",
   34895 => x"0c30c3",
   34896 => x"0c30c3",
   34897 => x"0c30c3",
   34898 => x"0c30c3",
   34899 => x"0c30c3",
   34900 => x"0c30c3",
   34901 => x"0c30c3",
   34902 => x"0c30c3",
   34903 => x"0c30c3",
   34904 => x"0c30c3",
   34905 => x"0c30c3",
   34906 => x"0c30c3",
   34907 => x"0c30c3",
   34908 => x"0c30c3",
   34909 => x"0c30c3",
   34910 => x"0c30c3",
   34911 => x"0c30c3",
   34912 => x"0c30c3",
   34913 => x"0c30c3",
   34914 => x"0c30c3",
   34915 => x"0c30c3",
   34916 => x"0c30c3",
   34917 => x"0c30c3",
   34918 => x"0c30c3",
   34919 => x"0c30c3",
   34920 => x"0c30c3",
   34921 => x"0c30c3",
   34922 => x"0c30c3",
   34923 => x"0c30c3",
   34924 => x"0c30c3",
   34925 => x"0c30c3",
   34926 => x"0c30c3",
   34927 => x"0c30c3",
   34928 => x"0c30c3",
   34929 => x"0c30c3",
   34930 => x"0c30c3",
   34931 => x"0c30c3",
   34932 => x"0c30c3",
   34933 => x"0c30c3",
   34934 => x"0c30c3",
   34935 => x"0c30c3",
   34936 => x"0d7fff",
   34937 => x"ffffff",
   34938 => x"ffffff",
   34939 => x"ffffff",
   34940 => x"ffffff",
   34941 => x"ffffff",
   34942 => x"ffffff",
   34943 => x"ffffff",
   34944 => x"ffffff",
   34945 => x"ffffff",
   34946 => x"ffffff",
   34947 => x"ffffff",
   34948 => x"ffffff",
   34949 => x"fffa95",
   34950 => x"abffff",
   34951 => x"ffffff",
   34952 => x"ffffff",
   34953 => x"ffffff",
   34954 => x"ffffff",
   34955 => x"ffffff",
   34956 => x"ffffff",
   34957 => x"ffffff",
   34958 => x"ffffff",
   34959 => x"ffffff",
   34960 => x"ffffff",
   34961 => x"ffffff",
   34962 => x"ffffff",
   34963 => x"ffffff",
   34964 => x"ffffff",
   34965 => x"ffffff",
   34966 => x"ffffff",
   34967 => x"ffffff",
   34968 => x"ffffff",
   34969 => x"ffffff",
   34970 => x"ffffff",
   34971 => x"ffffff",
   34972 => x"ffffff",
   34973 => x"ffffff",
   34974 => x"ffffff",
   34975 => x"ffffff",
   34976 => x"ffffff",
   34977 => x"ffffff",
   34978 => x"ffffff",
   34979 => x"ffffff",
   34980 => x"ffffff",
   34981 => x"ffffff",
   34982 => x"ffffff",
   34983 => x"ffffff",
   34984 => x"ffffff",
   34985 => x"ffffff",
   34986 => x"ffffff",
   34987 => x"ffffff",
   34988 => x"ffffff",
   34989 => x"ffffff",
   34990 => x"ffffff",
   34991 => x"ffffff",
   34992 => x"ffffff",
   34993 => x"ffffff",
   34994 => x"ffffff",
   34995 => x"ffffff",
   34996 => x"ffffff",
   34997 => x"ffffff",
   34998 => x"ffffff",
   34999 => x"ffffff",
   35000 => x"ffffff",
   35001 => x"ffffff",
   35002 => x"ffffff",
   35003 => x"ffffff",
   35004 => x"ffffff",
   35005 => x"ffffff",
   35006 => x"ffffff",
   35007 => x"ffffff",
   35008 => x"ffffff",
   35009 => x"ffffff",
   35010 => x"ffffff",
   35011 => x"ffffff",
   35012 => x"ffffff",
   35013 => x"ffffff",
   35014 => x"ffffff",
   35015 => x"ffffff",
   35016 => x"ffffff",
   35017 => x"ffffff",
   35018 => x"ffffff",
   35019 => x"ffffff",
   35020 => x"ffffff",
   35021 => x"ffffff",
   35022 => x"ffffff",
   35023 => x"ffffff",
   35024 => x"ffffff",
   35025 => x"ffffff",
   35026 => x"ffffff",
   35027 => x"ffffff",
   35028 => x"ffffff",
   35029 => x"ffffff",
   35030 => x"ffffff",
   35031 => x"ffffff",
   35032 => x"ffffff",
   35033 => x"ffffff",
   35034 => x"ffffff",
   35035 => x"ffffff",
   35036 => x"ffffff",
   35037 => x"ffffff",
   35038 => x"ffffff",
   35039 => x"ffffff",
   35040 => x"ffffff",
   35041 => x"ffffff",
   35042 => x"ffffff",
   35043 => x"ffffff",
   35044 => x"ffffff",
   35045 => x"ffffff",
   35046 => x"ffffff",
   35047 => x"ffffff",
   35048 => x"ffffff",
   35049 => x"ffffff",
   35050 => x"ffffff",
   35051 => x"ffffff",
   35052 => x"fd70c3",
   35053 => x"0c30c3",
   35054 => x"0c30c3",
   35055 => x"0c30c3",
   35056 => x"0c30c3",
   35057 => x"0c30c3",
   35058 => x"0c30c3",
   35059 => x"0c30c3",
   35060 => x"0c30c3",
   35061 => x"0c30c3",
   35062 => x"0c30c3",
   35063 => x"0c30c3",
   35064 => x"0c30c3",
   35065 => x"0c30c3",
   35066 => x"0c30c3",
   35067 => x"0c30c3",
   35068 => x"0c30c3",
   35069 => x"0c30c3",
   35070 => x"0c30c3",
   35071 => x"0c30c3",
   35072 => x"0c30c3",
   35073 => x"0c30c3",
   35074 => x"0c30c3",
   35075 => x"0c30c3",
   35076 => x"0c30c3",
   35077 => x"0c30c3",
   35078 => x"0c30c3",
   35079 => x"0c30c3",
   35080 => x"0c30c3",
   35081 => x"0c30c3",
   35082 => x"0c30c3",
   35083 => x"0c30c3",
   35084 => x"0c30c3",
   35085 => x"0c30c3",
   35086 => x"0c30c3",
   35087 => x"0c30c3",
   35088 => x"0c30c3",
   35089 => x"0c30c3",
   35090 => x"0c30c3",
   35091 => x"0c30c3",
   35092 => x"0c30c3",
   35093 => x"0c30c3",
   35094 => x"0c30c3",
   35095 => x"0c30c3",
   35096 => x"0ebfff",
   35097 => x"ffffff",
   35098 => x"ffffff",
   35099 => x"ffffff",
   35100 => x"ffffff",
   35101 => x"ffffff",
   35102 => x"ffffff",
   35103 => x"ffffff",
   35104 => x"ffffff",
   35105 => x"ffffff",
   35106 => x"ffffff",
   35107 => x"ffffff",
   35108 => x"ffffff",
   35109 => x"fffa95",
   35110 => x"abffff",
   35111 => x"ffffff",
   35112 => x"ffffff",
   35113 => x"ffffff",
   35114 => x"ffffff",
   35115 => x"ffffff",
   35116 => x"ffffff",
   35117 => x"ffffff",
   35118 => x"ffffff",
   35119 => x"ffffff",
   35120 => x"ffffff",
   35121 => x"ffffee",
   35122 => x"75d75d",
   35123 => x"75d75d",
   35124 => x"75d75d",
   35125 => x"75d75d",
   35126 => x"75d75d",
   35127 => x"75d75d",
   35128 => x"75d75d",
   35129 => x"75d75d",
   35130 => x"75d75d",
   35131 => x"75d75d",
   35132 => x"75d75d",
   35133 => x"75d75d",
   35134 => x"75d75d",
   35135 => x"75d75d",
   35136 => x"75d75d",
   35137 => x"75d75d",
   35138 => x"75d75d",
   35139 => x"75d75d",
   35140 => x"75d75d",
   35141 => x"75d75d",
   35142 => x"75d75d",
   35143 => x"75d659",
   35144 => x"659659",
   35145 => x"659659",
   35146 => x"659659",
   35147 => x"659659",
   35148 => x"659659",
   35149 => x"659659",
   35150 => x"659659",
   35151 => x"659659",
   35152 => x"659659",
   35153 => x"659659",
   35154 => x"659659",
   35155 => x"659659",
   35156 => x"659659",
   35157 => x"659659",
   35158 => x"659659",
   35159 => x"659659",
   35160 => x"659659",
   35161 => x"659659",
   35162 => x"659659",
   35163 => x"659659",
   35164 => x"659659",
   35165 => x"659659",
   35166 => x"659659",
   35167 => x"659659",
   35168 => x"659659",
   35169 => x"659659",
   35170 => x"659659",
   35171 => x"659659",
   35172 => x"659659",
   35173 => x"659659",
   35174 => x"659659",
   35175 => x"659659",
   35176 => x"659659",
   35177 => x"659659",
   35178 => x"659659",
   35179 => x"659659",
   35180 => x"659659",
   35181 => x"659659",
   35182 => x"659659",
   35183 => x"659659",
   35184 => x"659659",
   35185 => x"659659",
   35186 => x"659659",
   35187 => x"659659",
   35188 => x"659555",
   35189 => x"555abf",
   35190 => x"ffffff",
   35191 => x"ffffff",
   35192 => x"ffffff",
   35193 => x"ffffff",
   35194 => x"ffffff",
   35195 => x"ffffff",
   35196 => x"ffffff",
   35197 => x"ffffff",
   35198 => x"ffffff",
   35199 => x"ffffff",
   35200 => x"ffffff",
   35201 => x"ffffff",
   35202 => x"ffffff",
   35203 => x"ffffff",
   35204 => x"ffffff",
   35205 => x"ffffff",
   35206 => x"ffffff",
   35207 => x"ffffff",
   35208 => x"ffffff",
   35209 => x"ffffff",
   35210 => x"ffffff",
   35211 => x"ffffff",
   35212 => x"fd70c3",
   35213 => x"0c30c3",
   35214 => x"0c30c3",
   35215 => x"0c30c3",
   35216 => x"0c30c3",
   35217 => x"0c30c3",
   35218 => x"0c30c3",
   35219 => x"0c30c3",
   35220 => x"0c30c3",
   35221 => x"0c30c3",
   35222 => x"0c30c3",
   35223 => x"0c30c3",
   35224 => x"0c30c3",
   35225 => x"0c30c3",
   35226 => x"0c30c3",
   35227 => x"0c30c3",
   35228 => x"0c30c3",
   35229 => x"0c30c3",
   35230 => x"0c30c3",
   35231 => x"0c30c3",
   35232 => x"0c30c3",
   35233 => x"0c30c3",
   35234 => x"0c30c3",
   35235 => x"0c30c3",
   35236 => x"0c30c3",
   35237 => x"0c30c3",
   35238 => x"0c30c3",
   35239 => x"0c30c3",
   35240 => x"0c30c3",
   35241 => x"0c30c3",
   35242 => x"0c30c3",
   35243 => x"0c30c3",
   35244 => x"0c30c3",
   35245 => x"0c30c3",
   35246 => x"0c30c3",
   35247 => x"0c30c3",
   35248 => x"0c30c3",
   35249 => x"0c30c3",
   35250 => x"0c30c3",
   35251 => x"0c30c3",
   35252 => x"0c30c3",
   35253 => x"0c30c3",
   35254 => x"0c30c3",
   35255 => x"0c30c3",
   35256 => x"0ebfff",
   35257 => x"ffffff",
   35258 => x"ffffff",
   35259 => x"ffffff",
   35260 => x"ffffff",
   35261 => x"ffffff",
   35262 => x"ffffff",
   35263 => x"ffffff",
   35264 => x"ffffff",
   35265 => x"ffffff",
   35266 => x"ffffff",
   35267 => x"ffffff",
   35268 => x"ffffff",
   35269 => x"fffa95",
   35270 => x"abffff",
   35271 => x"ffffff",
   35272 => x"ffffff",
   35273 => x"ffffff",
   35274 => x"ffffff",
   35275 => x"ffffff",
   35276 => x"ffffff",
   35277 => x"ffffff",
   35278 => x"ffffff",
   35279 => x"ffffff",
   35280 => x"ffffff",
   35281 => x"fffb9d",
   35282 => x"30c30c",
   35283 => x"30c30c",
   35284 => x"30c30c",
   35285 => x"30c30c",
   35286 => x"30c30c",
   35287 => x"30c30c",
   35288 => x"30c30c",
   35289 => x"30c30c",
   35290 => x"30c30c",
   35291 => x"30c30c",
   35292 => x"30c30c",
   35293 => x"30c308",
   35294 => x"208208",
   35295 => x"208208",
   35296 => x"208208",
   35297 => x"208208",
   35298 => x"208208",
   35299 => x"208208",
   35300 => x"208208",
   35301 => x"208208",
   35302 => x"208208",
   35303 => x"208208",
   35304 => x"208208",
   35305 => x"208208",
   35306 => x"208208",
   35307 => x"208208",
   35308 => x"208208",
   35309 => x"208208",
   35310 => x"208208",
   35311 => x"208208",
   35312 => x"208208",
   35313 => x"208208",
   35314 => x"208208",
   35315 => x"208208",
   35316 => x"208208",
   35317 => x"208208",
   35318 => x"104104",
   35319 => x"104104",
   35320 => x"104104",
   35321 => x"104104",
   35322 => x"104104",
   35323 => x"104104",
   35324 => x"104104",
   35325 => x"104104",
   35326 => x"104104",
   35327 => x"104104",
   35328 => x"104104",
   35329 => x"104104",
   35330 => x"104104",
   35331 => x"104104",
   35332 => x"104104",
   35333 => x"104104",
   35334 => x"104104",
   35335 => x"104104",
   35336 => x"104104",
   35337 => x"104104",
   35338 => x"104104",
   35339 => x"104104",
   35340 => x"104104",
   35341 => x"104104",
   35342 => x"000000",
   35343 => x"000000",
   35344 => x"000000",
   35345 => x"000000",
   35346 => x"000000",
   35347 => x"000000",
   35348 => x"000000",
   35349 => x"000abf",
   35350 => x"ffffff",
   35351 => x"ffffff",
   35352 => x"ffffff",
   35353 => x"ffffff",
   35354 => x"ffffff",
   35355 => x"ffffff",
   35356 => x"ffffff",
   35357 => x"ffffff",
   35358 => x"ffffff",
   35359 => x"ffffff",
   35360 => x"ffffff",
   35361 => x"ffffff",
   35362 => x"ffffff",
   35363 => x"ffffff",
   35364 => x"ffffff",
   35365 => x"ffffff",
   35366 => x"ffffff",
   35367 => x"ffffff",
   35368 => x"ffffff",
   35369 => x"ffffff",
   35370 => x"ffffff",
   35371 => x"ffffff",
   35372 => x"feb0c3",
   35373 => x"0c30c3",
   35374 => x"0c30c3",
   35375 => x"0c30c3",
   35376 => x"0c30c3",
   35377 => x"0c30c3",
   35378 => x"0c30c3",
   35379 => x"0c30c3",
   35380 => x"0c30c3",
   35381 => x"0c30c3",
   35382 => x"0c30c3",
   35383 => x"0c30c3",
   35384 => x"0c30c3",
   35385 => x"0c30c3",
   35386 => x"0c30c3",
   35387 => x"0c30c3",
   35388 => x"0c30c3",
   35389 => x"0c30c3",
   35390 => x"0c30c3",
   35391 => x"0c30c3",
   35392 => x"0c30c3",
   35393 => x"0c30c3",
   35394 => x"0c30c3",
   35395 => x"0c30c3",
   35396 => x"0c30c3",
   35397 => x"0c30c3",
   35398 => x"0c30c3",
   35399 => x"0c30c3",
   35400 => x"0c30c3",
   35401 => x"0c30c3",
   35402 => x"0c30c3",
   35403 => x"0c30c3",
   35404 => x"0c30c3",
   35405 => x"0c30c3",
   35406 => x"0c30c3",
   35407 => x"0c30c3",
   35408 => x"0c30c3",
   35409 => x"0c30c3",
   35410 => x"0c30c3",
   35411 => x"0c30c3",
   35412 => x"0c30c3",
   35413 => x"0c30c3",
   35414 => x"0c30c3",
   35415 => x"0c30c3",
   35416 => x"5fffff",
   35417 => x"ffffff",
   35418 => x"ffffff",
   35419 => x"ffffff",
   35420 => x"ffffff",
   35421 => x"ffffff",
   35422 => x"ffffff",
   35423 => x"ffffff",
   35424 => x"ffffff",
   35425 => x"ffffff",
   35426 => x"ffffff",
   35427 => x"ffffff",
   35428 => x"ffffff",
   35429 => x"fffa95",
   35430 => x"abffff",
   35431 => x"ffffff",
   35432 => x"ffffff",
   35433 => x"ffffff",
   35434 => x"ffffff",
   35435 => x"ffffff",
   35436 => x"ffffff",
   35437 => x"ffffff",
   35438 => x"ffffff",
   35439 => x"ffffff",
   35440 => x"ffffff",
   35441 => x"fffb8c",
   35442 => x"30c30c",
   35443 => x"30c30c",
   35444 => x"30c30c",
   35445 => x"30c30c",
   35446 => x"30c30c",
   35447 => x"30c30c",
   35448 => x"30c30c",
   35449 => x"30c30c",
   35450 => x"30c30c",
   35451 => x"30c30c",
   35452 => x"30c30c",
   35453 => x"208208",
   35454 => x"208208",
   35455 => x"208208",
   35456 => x"208208",
   35457 => x"208208",
   35458 => x"208208",
   35459 => x"208208",
   35460 => x"208208",
   35461 => x"208208",
   35462 => x"208208",
   35463 => x"208208",
   35464 => x"208208",
   35465 => x"208208",
   35466 => x"208208",
   35467 => x"208208",
   35468 => x"208208",
   35469 => x"208208",
   35470 => x"208208",
   35471 => x"208208",
   35472 => x"208208",
   35473 => x"208208",
   35474 => x"208208",
   35475 => x"208104",
   35476 => x"104104",
   35477 => x"104104",
   35478 => x"104104",
   35479 => x"104104",
   35480 => x"104104",
   35481 => x"104104",
   35482 => x"104104",
   35483 => x"104104",
   35484 => x"104104",
   35485 => x"104104",
   35486 => x"104104",
   35487 => x"104104",
   35488 => x"104104",
   35489 => x"104104",
   35490 => x"104104",
   35491 => x"104104",
   35492 => x"104104",
   35493 => x"104104",
   35494 => x"104104",
   35495 => x"104104",
   35496 => x"104104",
   35497 => x"104104",
   35498 => x"104000",
   35499 => x"000000",
   35500 => x"000000",
   35501 => x"000000",
   35502 => x"000000",
   35503 => x"000000",
   35504 => x"000000",
   35505 => x"000000",
   35506 => x"000000",
   35507 => x"000000",
   35508 => x"000000",
   35509 => x"00057f",
   35510 => x"ffffff",
   35511 => x"ffffff",
   35512 => x"ffffff",
   35513 => x"ffffff",
   35514 => x"ffffff",
   35515 => x"ffffff",
   35516 => x"ffffff",
   35517 => x"ffffff",
   35518 => x"ffffff",
   35519 => x"ffffff",
   35520 => x"ffffff",
   35521 => x"ffffff",
   35522 => x"ffffff",
   35523 => x"ffffff",
   35524 => x"ffffff",
   35525 => x"ffffff",
   35526 => x"ffffff",
   35527 => x"ffffff",
   35528 => x"ffffff",
   35529 => x"ffffff",
   35530 => x"ffffff",
   35531 => x"ffffff",
   35532 => x"fff5c3",
   35533 => x"0c30c3",
   35534 => x"0c30c3",
   35535 => x"0c30c3",
   35536 => x"0c30c3",
   35537 => x"0c30c3",
   35538 => x"0c30c3",
   35539 => x"0c30c3",
   35540 => x"0c30c3",
   35541 => x"0c30c3",
   35542 => x"0c30c3",
   35543 => x"0c30c3",
   35544 => x"0c30c3",
   35545 => x"0c30c3",
   35546 => x"0c30c3",
   35547 => x"0c30c3",
   35548 => x"0c30c3",
   35549 => x"0c30c3",
   35550 => x"0c30c3",
   35551 => x"0c30c3",
   35552 => x"0c30c3",
   35553 => x"0c30c3",
   35554 => x"0c30c3",
   35555 => x"0c30c3",
   35556 => x"0c30c3",
   35557 => x"0c30c3",
   35558 => x"0c30c3",
   35559 => x"0c30c3",
   35560 => x"0c30c3",
   35561 => x"0c30c3",
   35562 => x"0c30c3",
   35563 => x"0c30c3",
   35564 => x"0c30c3",
   35565 => x"0c30c3",
   35566 => x"0c30c3",
   35567 => x"0c30c3",
   35568 => x"0c30c3",
   35569 => x"0c30c3",
   35570 => x"0c30c3",
   35571 => x"0c30c3",
   35572 => x"0c30c3",
   35573 => x"0c30c3",
   35574 => x"0c30c3",
   35575 => x"0c30c3",
   35576 => x"afffff",
   35577 => x"ffffff",
   35578 => x"ffffff",
   35579 => x"ffffff",
   35580 => x"ffffff",
   35581 => x"ffffff",
   35582 => x"ffffff",
   35583 => x"ffffff",
   35584 => x"ffffff",
   35585 => x"ffffff",
   35586 => x"ffffff",
   35587 => x"ffffff",
   35588 => x"ffffff",
   35589 => x"fffa95",
   35590 => x"abffff",
   35591 => x"ffffff",
   35592 => x"ffffff",
   35593 => x"ffffff",
   35594 => x"ffffff",
   35595 => x"ffffff",
   35596 => x"ffffff",
   35597 => x"ffffff",
   35598 => x"ffffff",
   35599 => x"ffffff",
   35600 => x"ffffff",
   35601 => x"fffb8c",
   35602 => x"30c30c",
   35603 => x"30c30c",
   35604 => x"30c30c",
   35605 => x"30c30c",
   35606 => x"30c30c",
   35607 => x"30c30c",
   35608 => x"30c30c",
   35609 => x"30c30c",
   35610 => x"30c30c",
   35611 => x"30c30c",
   35612 => x"30c30c",
   35613 => x"208208",
   35614 => x"208208",
   35615 => x"208208",
   35616 => x"208208",
   35617 => x"208208",
   35618 => x"208208",
   35619 => x"208208",
   35620 => x"208208",
   35621 => x"208208",
   35622 => x"208208",
   35623 => x"208208",
   35624 => x"208208",
   35625 => x"208208",
   35626 => x"208208",
   35627 => x"208208",
   35628 => x"208208",
   35629 => x"208208",
   35630 => x"208208",
   35631 => x"208208",
   35632 => x"208208",
   35633 => x"208208",
   35634 => x"208208",
   35635 => x"208104",
   35636 => x"104104",
   35637 => x"104104",
   35638 => x"104104",
   35639 => x"104104",
   35640 => x"104104",
   35641 => x"104104",
   35642 => x"104104",
   35643 => x"104104",
   35644 => x"104104",
   35645 => x"104104",
   35646 => x"104104",
   35647 => x"104104",
   35648 => x"104104",
   35649 => x"104104",
   35650 => x"104104",
   35651 => x"104104",
   35652 => x"104104",
   35653 => x"104104",
   35654 => x"104104",
   35655 => x"104104",
   35656 => x"104104",
   35657 => x"104104",
   35658 => x"104000",
   35659 => x"000000",
   35660 => x"000000",
   35661 => x"000000",
   35662 => x"000000",
   35663 => x"000000",
   35664 => x"000000",
   35665 => x"000000",
   35666 => x"000000",
   35667 => x"000000",
   35668 => x"000000",
   35669 => x"00057f",
   35670 => x"ffffff",
   35671 => x"ffffff",
   35672 => x"ffffff",
   35673 => x"ffffff",
   35674 => x"ffffff",
   35675 => x"ffffff",
   35676 => x"ffffff",
   35677 => x"ffffff",
   35678 => x"ffffff",
   35679 => x"ffffff",
   35680 => x"ffffff",
   35681 => x"ffffff",
   35682 => x"ffffff",
   35683 => x"ffffff",
   35684 => x"ffffff",
   35685 => x"ffffff",
   35686 => x"ffffff",
   35687 => x"ffffff",
   35688 => x"ffffff",
   35689 => x"ffffff",
   35690 => x"ffffff",
   35691 => x"ffffff",
   35692 => x"fffac3",
   35693 => x"0c30c3",
   35694 => x"0c30c3",
   35695 => x"0c30c3",
   35696 => x"0c30c3",
   35697 => x"0c30c3",
   35698 => x"0c30c3",
   35699 => x"0c30c3",
   35700 => x"0c30c3",
   35701 => x"0c30c3",
   35702 => x"0c30c3",
   35703 => x"0c30c3",
   35704 => x"0c30c3",
   35705 => x"0c30c3",
   35706 => x"0c30c3",
   35707 => x"0c30c3",
   35708 => x"0c30c3",
   35709 => x"0c30c3",
   35710 => x"0c30c3",
   35711 => x"0c30c3",
   35712 => x"0c30c3",
   35713 => x"0c30c3",
   35714 => x"0c30c3",
   35715 => x"0c30c3",
   35716 => x"0c30c3",
   35717 => x"0c30c3",
   35718 => x"0c30c3",
   35719 => x"0c30c3",
   35720 => x"0c30c3",
   35721 => x"0c30c3",
   35722 => x"0c30c3",
   35723 => x"0c30c3",
   35724 => x"0c30c3",
   35725 => x"0c30c3",
   35726 => x"0c30c3",
   35727 => x"0c30c3",
   35728 => x"0c30c3",
   35729 => x"0c30c3",
   35730 => x"0c30c3",
   35731 => x"0c30c3",
   35732 => x"0c30c3",
   35733 => x"0c30c3",
   35734 => x"0c30c3",
   35735 => x"0c30d7",
   35736 => x"afffff",
   35737 => x"ffffff",
   35738 => x"ffffff",
   35739 => x"ffffff",
   35740 => x"ffffff",
   35741 => x"ffffff",
   35742 => x"ffffff",
   35743 => x"ffffff",
   35744 => x"ffffff",
   35745 => x"ffffff",
   35746 => x"ffffff",
   35747 => x"ffffff",
   35748 => x"ffffff",
   35749 => x"fffa95",
   35750 => x"abffff",
   35751 => x"ffffff",
   35752 => x"ffffff",
   35753 => x"ffffff",
   35754 => x"ffffff",
   35755 => x"ffffff",
   35756 => x"ffffff",
   35757 => x"ffffff",
   35758 => x"ffffff",
   35759 => x"ffffff",
   35760 => x"ffffff",
   35761 => x"fffb8c",
   35762 => x"30c30c",
   35763 => x"30c30c",
   35764 => x"30c30c",
   35765 => x"30c30c",
   35766 => x"30c30c",
   35767 => x"30c30c",
   35768 => x"30c30c",
   35769 => x"30c30c",
   35770 => x"30c30c",
   35771 => x"30c30c",
   35772 => x"30c30c",
   35773 => x"208208",
   35774 => x"208208",
   35775 => x"208208",
   35776 => x"208208",
   35777 => x"208208",
   35778 => x"208208",
   35779 => x"208208",
   35780 => x"208208",
   35781 => x"208208",
   35782 => x"208208",
   35783 => x"208208",
   35784 => x"208208",
   35785 => x"208208",
   35786 => x"208208",
   35787 => x"208208",
   35788 => x"208208",
   35789 => x"208208",
   35790 => x"208208",
   35791 => x"208208",
   35792 => x"208208",
   35793 => x"208208",
   35794 => x"208208",
   35795 => x"208104",
   35796 => x"104104",
   35797 => x"104104",
   35798 => x"104104",
   35799 => x"104104",
   35800 => x"104104",
   35801 => x"104104",
   35802 => x"104104",
   35803 => x"104104",
   35804 => x"104104",
   35805 => x"104104",
   35806 => x"104104",
   35807 => x"104104",
   35808 => x"104104",
   35809 => x"104104",
   35810 => x"104104",
   35811 => x"104104",
   35812 => x"104104",
   35813 => x"104104",
   35814 => x"104104",
   35815 => x"104104",
   35816 => x"104104",
   35817 => x"104104",
   35818 => x"104000",
   35819 => x"000000",
   35820 => x"000000",
   35821 => x"000000",
   35822 => x"000000",
   35823 => x"000000",
   35824 => x"000000",
   35825 => x"000000",
   35826 => x"000000",
   35827 => x"000000",
   35828 => x"000000",
   35829 => x"00057f",
   35830 => x"ffffff",
   35831 => x"ffffff",
   35832 => x"ffffff",
   35833 => x"ffffff",
   35834 => x"ffffff",
   35835 => x"ffffff",
   35836 => x"ffffff",
   35837 => x"ffffff",
   35838 => x"ffffff",
   35839 => x"ffffff",
   35840 => x"ffffff",
   35841 => x"ffffff",
   35842 => x"ffffff",
   35843 => x"ffffff",
   35844 => x"ffffff",
   35845 => x"ffffff",
   35846 => x"ffffff",
   35847 => x"ffffff",
   35848 => x"ffffff",
   35849 => x"ffffff",
   35850 => x"ffffff",
   35851 => x"ffffff",
   35852 => x"fffac3",
   35853 => x"0c30c3",
   35854 => x"0c30c3",
   35855 => x"0c30c3",
   35856 => x"0c30c3",
   35857 => x"0c30c3",
   35858 => x"0c30c3",
   35859 => x"0c30c3",
   35860 => x"0c30c3",
   35861 => x"0c30c3",
   35862 => x"0c30c3",
   35863 => x"0c30c3",
   35864 => x"0c30c3",
   35865 => x"0c30c3",
   35866 => x"0c30c3",
   35867 => x"0c30c3",
   35868 => x"0c30c3",
   35869 => x"0c30c3",
   35870 => x"0c30c3",
   35871 => x"0c30c3",
   35872 => x"0c30c3",
   35873 => x"0c30c3",
   35874 => x"0c30c3",
   35875 => x"0c30c3",
   35876 => x"0c30c3",
   35877 => x"0c30c3",
   35878 => x"0c30c3",
   35879 => x"0c30c3",
   35880 => x"0c30c3",
   35881 => x"0c30c3",
   35882 => x"0c30c3",
   35883 => x"0c30c3",
   35884 => x"0c30c3",
   35885 => x"0c30c3",
   35886 => x"0c30c3",
   35887 => x"0c30c3",
   35888 => x"0c30c3",
   35889 => x"0c30c3",
   35890 => x"0c30c3",
   35891 => x"0c30c3",
   35892 => x"0c30c3",
   35893 => x"0c30c3",
   35894 => x"0c30c3",
   35895 => x"0c30d7",
   35896 => x"ffffff",
   35897 => x"ffffff",
   35898 => x"ffffff",
   35899 => x"ffffff",
   35900 => x"ffffff",
   35901 => x"ffffff",
   35902 => x"ffffff",
   35903 => x"ffffff",
   35904 => x"ffffff",
   35905 => x"ffffff",
   35906 => x"ffffff",
   35907 => x"ffffff",
   35908 => x"ffffff",
   35909 => x"fffa95",
   35910 => x"abffff",
   35911 => x"ffffff",
   35912 => x"ffffff",
   35913 => x"ffffff",
   35914 => x"ffffff",
   35915 => x"ffffff",
   35916 => x"ffffff",
   35917 => x"ffffff",
   35918 => x"ffffff",
   35919 => x"ffffff",
   35920 => x"ffffff",
   35921 => x"fffb8c",
   35922 => x"30c30c",
   35923 => x"30c30c",
   35924 => x"30c30c",
   35925 => x"30c30c",
   35926 => x"30c30c",
   35927 => x"30c30c",
   35928 => x"30c30c",
   35929 => x"30c30c",
   35930 => x"30c30c",
   35931 => x"30c30c",
   35932 => x"30c30c",
   35933 => x"208208",
   35934 => x"208208",
   35935 => x"208208",
   35936 => x"208208",
   35937 => x"208208",
   35938 => x"208208",
   35939 => x"208208",
   35940 => x"208208",
   35941 => x"208208",
   35942 => x"208208",
   35943 => x"208208",
   35944 => x"208208",
   35945 => x"208208",
   35946 => x"208208",
   35947 => x"208208",
   35948 => x"208208",
   35949 => x"208208",
   35950 => x"208208",
   35951 => x"208208",
   35952 => x"208208",
   35953 => x"208208",
   35954 => x"208208",
   35955 => x"208104",
   35956 => x"104104",
   35957 => x"104104",
   35958 => x"104104",
   35959 => x"104104",
   35960 => x"104104",
   35961 => x"104104",
   35962 => x"104104",
   35963 => x"104104",
   35964 => x"104104",
   35965 => x"104104",
   35966 => x"104104",
   35967 => x"104104",
   35968 => x"104104",
   35969 => x"104104",
   35970 => x"104104",
   35971 => x"104104",
   35972 => x"104104",
   35973 => x"104104",
   35974 => x"104104",
   35975 => x"104104",
   35976 => x"104104",
   35977 => x"104104",
   35978 => x"104000",
   35979 => x"000000",
   35980 => x"000000",
   35981 => x"000000",
   35982 => x"000000",
   35983 => x"000000",
   35984 => x"000000",
   35985 => x"000000",
   35986 => x"000000",
   35987 => x"000000",
   35988 => x"000000",
   35989 => x"00057f",
   35990 => x"ffffff",
   35991 => x"ffffff",
   35992 => x"ffffff",
   35993 => x"ffffff",
   35994 => x"ffffff",
   35995 => x"ffffff",
   35996 => x"ffffff",
   35997 => x"ffffff",
   35998 => x"ffffff",
   35999 => x"ffffff",
   36000 => x"ffffff",
   36001 => x"ffffff",
   36002 => x"ffffff",
   36003 => x"ffffff",
   36004 => x"ffffff",
   36005 => x"ffffff",
   36006 => x"ffffff",
   36007 => x"ffffff",
   36008 => x"ffffff",
   36009 => x"ffffff",
   36010 => x"ffffff",
   36011 => x"ffffff",
   36012 => x"ffffd7",
   36013 => x"0c30c3",
   36014 => x"0c30c3",
   36015 => x"0c30c3",
   36016 => x"0c30c3",
   36017 => x"0c30c3",
   36018 => x"0c30c3",
   36019 => x"0c30c3",
   36020 => x"0c30c3",
   36021 => x"0c30c3",
   36022 => x"0c30c3",
   36023 => x"0c30c3",
   36024 => x"0c30c3",
   36025 => x"0c30c3",
   36026 => x"0c30c3",
   36027 => x"0c30c3",
   36028 => x"0c30c3",
   36029 => x"0c30c3",
   36030 => x"0c30c3",
   36031 => x"0c30c3",
   36032 => x"0c30c3",
   36033 => x"0c30c3",
   36034 => x"0c30c3",
   36035 => x"0c30c3",
   36036 => x"0c30c3",
   36037 => x"0c30c3",
   36038 => x"0c30c3",
   36039 => x"0c30c3",
   36040 => x"0c30c3",
   36041 => x"0c30c3",
   36042 => x"0c30c3",
   36043 => x"0c30c3",
   36044 => x"0c30c3",
   36045 => x"0c30c3",
   36046 => x"0c30c3",
   36047 => x"0c30c3",
   36048 => x"0c30c3",
   36049 => x"0c30c3",
   36050 => x"0c30c3",
   36051 => x"0c30c3",
   36052 => x"0c30c3",
   36053 => x"0c30c3",
   36054 => x"0c30c3",
   36055 => x"0c30eb",
   36056 => x"ffffff",
   36057 => x"ffffff",
   36058 => x"ffffff",
   36059 => x"ffffff",
   36060 => x"ffffff",
   36061 => x"ffffff",
   36062 => x"ffffff",
   36063 => x"ffffff",
   36064 => x"ffffff",
   36065 => x"ffffff",
   36066 => x"ffffff",
   36067 => x"ffffff",
   36068 => x"ffffff",
   36069 => x"fffa95",
   36070 => x"abffff",
   36071 => x"ffffff",
   36072 => x"ffffff",
   36073 => x"ffffff",
   36074 => x"ffffff",
   36075 => x"ffffff",
   36076 => x"ffffff",
   36077 => x"ffffff",
   36078 => x"ffffff",
   36079 => x"ffffff",
   36080 => x"ffffff",
   36081 => x"fffb8c",
   36082 => x"30c30c",
   36083 => x"30c30c",
   36084 => x"30c30c",
   36085 => x"30c30c",
   36086 => x"30c30c",
   36087 => x"30c30c",
   36088 => x"30c30c",
   36089 => x"30c30c",
   36090 => x"30c30c",
   36091 => x"30c30c",
   36092 => x"30c30c",
   36093 => x"208208",
   36094 => x"208208",
   36095 => x"208208",
   36096 => x"208208",
   36097 => x"208208",
   36098 => x"208208",
   36099 => x"208208",
   36100 => x"208208",
   36101 => x"208208",
   36102 => x"208208",
   36103 => x"208208",
   36104 => x"208208",
   36105 => x"208208",
   36106 => x"208208",
   36107 => x"208208",
   36108 => x"208208",
   36109 => x"208208",
   36110 => x"208208",
   36111 => x"208208",
   36112 => x"208208",
   36113 => x"208208",
   36114 => x"208208",
   36115 => x"208104",
   36116 => x"104104",
   36117 => x"104104",
   36118 => x"104104",
   36119 => x"104104",
   36120 => x"104104",
   36121 => x"104104",
   36122 => x"104104",
   36123 => x"104104",
   36124 => x"104104",
   36125 => x"104104",
   36126 => x"104104",
   36127 => x"104104",
   36128 => x"104104",
   36129 => x"104104",
   36130 => x"104104",
   36131 => x"104104",
   36132 => x"104104",
   36133 => x"104104",
   36134 => x"104104",
   36135 => x"104104",
   36136 => x"104104",
   36137 => x"104104",
   36138 => x"104000",
   36139 => x"000000",
   36140 => x"000000",
   36141 => x"000000",
   36142 => x"000000",
   36143 => x"000000",
   36144 => x"000000",
   36145 => x"000000",
   36146 => x"000000",
   36147 => x"000000",
   36148 => x"000000",
   36149 => x"00057f",
   36150 => x"ffffff",
   36151 => x"ffffff",
   36152 => x"ffffff",
   36153 => x"ffffff",
   36154 => x"ffffff",
   36155 => x"ffffff",
   36156 => x"ffffff",
   36157 => x"ffffff",
   36158 => x"ffffff",
   36159 => x"ffffff",
   36160 => x"ffffff",
   36161 => x"ffffff",
   36162 => x"ffffff",
   36163 => x"ffffff",
   36164 => x"ffffff",
   36165 => x"ffffff",
   36166 => x"ffffff",
   36167 => x"ffffff",
   36168 => x"ffffff",
   36169 => x"ffffff",
   36170 => x"ffffff",
   36171 => x"ffffff",
   36172 => x"ffffeb",
   36173 => x"0c30c3",
   36174 => x"0c30c3",
   36175 => x"0c30c3",
   36176 => x"0c30c3",
   36177 => x"0c30c3",
   36178 => x"0c30c3",
   36179 => x"0c30c3",
   36180 => x"0c30c3",
   36181 => x"0c30c3",
   36182 => x"0c30c3",
   36183 => x"0c30c3",
   36184 => x"0c30c3",
   36185 => x"0c30c3",
   36186 => x"0c30c3",
   36187 => x"0c30c3",
   36188 => x"0c30c3",
   36189 => x"0c30c3",
   36190 => x"0c30c3",
   36191 => x"0c30c3",
   36192 => x"0c30c3",
   36193 => x"0c30c3",
   36194 => x"0c30c3",
   36195 => x"0c30c3",
   36196 => x"0c30c3",
   36197 => x"0c30c3",
   36198 => x"0c30c3",
   36199 => x"0c30c3",
   36200 => x"0c30c3",
   36201 => x"0c30c3",
   36202 => x"0c30c3",
   36203 => x"0c30c3",
   36204 => x"0c30c3",
   36205 => x"0c30c3",
   36206 => x"0c30c3",
   36207 => x"0c30c3",
   36208 => x"0c30c3",
   36209 => x"0c30c3",
   36210 => x"0c30c3",
   36211 => x"0c30c3",
   36212 => x"0c30c3",
   36213 => x"0c30c3",
   36214 => x"0c30c3",
   36215 => x"0c35eb",
   36216 => x"ffffff",
   36217 => x"ffffff",
   36218 => x"ffffff",
   36219 => x"ffffff",
   36220 => x"ffffff",
   36221 => x"ffffff",
   36222 => x"ffffff",
   36223 => x"ffffff",
   36224 => x"ffffff",
   36225 => x"ffffff",
   36226 => x"ffffff",
   36227 => x"ffffff",
   36228 => x"ffffff",
   36229 => x"fffa95",
   36230 => x"abffff",
   36231 => x"ffffff",
   36232 => x"ffffff",
   36233 => x"ffffff",
   36234 => x"ffffff",
   36235 => x"ffffff",
   36236 => x"ffffff",
   36237 => x"ffffff",
   36238 => x"ffffff",
   36239 => x"ffffff",
   36240 => x"ffffff",
   36241 => x"fffb8c",
   36242 => x"30c30c",
   36243 => x"30c30c",
   36244 => x"30c30c",
   36245 => x"30c30c",
   36246 => x"30c30c",
   36247 => x"30c30c",
   36248 => x"30c30c",
   36249 => x"30c30c",
   36250 => x"30c30c",
   36251 => x"30c30c",
   36252 => x"30c30c",
   36253 => x"208208",
   36254 => x"208208",
   36255 => x"208208",
   36256 => x"208208",
   36257 => x"208208",
   36258 => x"208208",
   36259 => x"208208",
   36260 => x"208208",
   36261 => x"208208",
   36262 => x"208208",
   36263 => x"208208",
   36264 => x"208208",
   36265 => x"208208",
   36266 => x"208208",
   36267 => x"208208",
   36268 => x"208208",
   36269 => x"208208",
   36270 => x"208208",
   36271 => x"208208",
   36272 => x"208208",
   36273 => x"208208",
   36274 => x"208208",
   36275 => x"208104",
   36276 => x"104104",
   36277 => x"104104",
   36278 => x"104104",
   36279 => x"104104",
   36280 => x"104104",
   36281 => x"104104",
   36282 => x"104104",
   36283 => x"104104",
   36284 => x"104104",
   36285 => x"104104",
   36286 => x"104104",
   36287 => x"104104",
   36288 => x"104104",
   36289 => x"104104",
   36290 => x"104104",
   36291 => x"104104",
   36292 => x"104104",
   36293 => x"104104",
   36294 => x"104104",
   36295 => x"104104",
   36296 => x"104104",
   36297 => x"104104",
   36298 => x"104000",
   36299 => x"000000",
   36300 => x"000000",
   36301 => x"000000",
   36302 => x"000000",
   36303 => x"000000",
   36304 => x"000000",
   36305 => x"000000",
   36306 => x"000000",
   36307 => x"000000",
   36308 => x"000000",
   36309 => x"00057f",
   36310 => x"ffffff",
   36311 => x"ffffff",
   36312 => x"ffffff",
   36313 => x"ffffff",
   36314 => x"ffffff",
   36315 => x"ffffff",
   36316 => x"ffffff",
   36317 => x"ffffff",
   36318 => x"ffffff",
   36319 => x"ffffff",
   36320 => x"ffffff",
   36321 => x"ffffff",
   36322 => x"ffffff",
   36323 => x"ffffff",
   36324 => x"ffffff",
   36325 => x"ffffff",
   36326 => x"ffffff",
   36327 => x"ffffff",
   36328 => x"ffffff",
   36329 => x"ffffff",
   36330 => x"ffffff",
   36331 => x"ffffff",
   36332 => x"ffffff",
   36333 => x"0c30c3",
   36334 => x"0c30c3",
   36335 => x"0c30c3",
   36336 => x"0c30c3",
   36337 => x"0c30c3",
   36338 => x"0c30c3",
   36339 => x"0c30c3",
   36340 => x"0c30c3",
   36341 => x"0c30c3",
   36342 => x"0c30c3",
   36343 => x"0c30c3",
   36344 => x"0c30c3",
   36345 => x"0c30c3",
   36346 => x"0c30c3",
   36347 => x"0c30c3",
   36348 => x"0c30c3",
   36349 => x"0c30c3",
   36350 => x"0c30c3",
   36351 => x"0c30c3",
   36352 => x"0c30c3",
   36353 => x"0c30c3",
   36354 => x"0c30c3",
   36355 => x"0c30c3",
   36356 => x"0c30c3",
   36357 => x"0c30c3",
   36358 => x"0c30c3",
   36359 => x"0c30c3",
   36360 => x"0c30c3",
   36361 => x"0c30c3",
   36362 => x"0c30c3",
   36363 => x"0c30c3",
   36364 => x"0c30c3",
   36365 => x"0c30c3",
   36366 => x"0c30c3",
   36367 => x"0c30c3",
   36368 => x"0c30c3",
   36369 => x"0c30c3",
   36370 => x"0c30c3",
   36371 => x"0c30c3",
   36372 => x"0c30c3",
   36373 => x"0c30c3",
   36374 => x"0c30c3",
   36375 => x"0c35ff",
   36376 => x"ffffff",
   36377 => x"ffffff",
   36378 => x"ffffff",
   36379 => x"ffffff",
   36380 => x"ffffff",
   36381 => x"ffffff",
   36382 => x"ffffff",
   36383 => x"ffffff",
   36384 => x"ffffff",
   36385 => x"ffffff",
   36386 => x"ffffff",
   36387 => x"ffffff",
   36388 => x"ffffff",
   36389 => x"fffa95",
   36390 => x"abffff",
   36391 => x"ffffff",
   36392 => x"ffffff",
   36393 => x"ffffff",
   36394 => x"ffffff",
   36395 => x"ffffff",
   36396 => x"ffffff",
   36397 => x"ffffff",
   36398 => x"ffffff",
   36399 => x"ffffff",
   36400 => x"ffffff",
   36401 => x"fffb8c",
   36402 => x"30c30c",
   36403 => x"30c30c",
   36404 => x"30c30c",
   36405 => x"30c30c",
   36406 => x"30c30c",
   36407 => x"30c30c",
   36408 => x"30c30c",
   36409 => x"30c30c",
   36410 => x"30c30c",
   36411 => x"30c30c",
   36412 => x"30c30c",
   36413 => x"208208",
   36414 => x"208208",
   36415 => x"208208",
   36416 => x"208208",
   36417 => x"208208",
   36418 => x"208208",
   36419 => x"208208",
   36420 => x"208208",
   36421 => x"208208",
   36422 => x"208208",
   36423 => x"208208",
   36424 => x"208208",
   36425 => x"208208",
   36426 => x"208208",
   36427 => x"208208",
   36428 => x"208208",
   36429 => x"208208",
   36430 => x"208208",
   36431 => x"208208",
   36432 => x"208208",
   36433 => x"208208",
   36434 => x"208208",
   36435 => x"208104",
   36436 => x"104104",
   36437 => x"104104",
   36438 => x"104104",
   36439 => x"104104",
   36440 => x"104104",
   36441 => x"104104",
   36442 => x"104104",
   36443 => x"104104",
   36444 => x"104104",
   36445 => x"104104",
   36446 => x"104104",
   36447 => x"104104",
   36448 => x"104104",
   36449 => x"104104",
   36450 => x"104104",
   36451 => x"104104",
   36452 => x"104104",
   36453 => x"104104",
   36454 => x"104104",
   36455 => x"104104",
   36456 => x"104104",
   36457 => x"104104",
   36458 => x"104000",
   36459 => x"000000",
   36460 => x"000000",
   36461 => x"000000",
   36462 => x"000000",
   36463 => x"000000",
   36464 => x"000000",
   36465 => x"000000",
   36466 => x"000000",
   36467 => x"000000",
   36468 => x"000000",
   36469 => x"00057f",
   36470 => x"ffffff",
   36471 => x"ffffff",
   36472 => x"ffffff",
   36473 => x"ffffff",
   36474 => x"ffffff",
   36475 => x"ffffff",
   36476 => x"ffffff",
   36477 => x"ffffff",
   36478 => x"ffffff",
   36479 => x"ffffff",
   36480 => x"ffffff",
   36481 => x"ffffff",
   36482 => x"ffffff",
   36483 => x"ffffff",
   36484 => x"ffffff",
   36485 => x"ffffff",
   36486 => x"ffffff",
   36487 => x"ffffff",
   36488 => x"ffffff",
   36489 => x"ffffff",
   36490 => x"ffffff",
   36491 => x"ffffff",
   36492 => x"ffffff",
   36493 => x"5c30c3",
   36494 => x"0c30c3",
   36495 => x"0c30c3",
   36496 => x"0c30c3",
   36497 => x"0c30c3",
   36498 => x"0c30c3",
   36499 => x"0c30c3",
   36500 => x"0c30c3",
   36501 => x"0c30c3",
   36502 => x"0c30c3",
   36503 => x"0c30c3",
   36504 => x"0c30c3",
   36505 => x"0c30c3",
   36506 => x"0c30c3",
   36507 => x"0c30c3",
   36508 => x"0c30c3",
   36509 => x"0c30c3",
   36510 => x"0c30c3",
   36511 => x"0c30c3",
   36512 => x"0c30c3",
   36513 => x"0c30c3",
   36514 => x"0c30c3",
   36515 => x"0c30c3",
   36516 => x"0c30c3",
   36517 => x"0c30c3",
   36518 => x"0c30c3",
   36519 => x"0c30c3",
   36520 => x"0c30c3",
   36521 => x"0c30c3",
   36522 => x"0c30c3",
   36523 => x"0c30c3",
   36524 => x"0c30c3",
   36525 => x"0c30c3",
   36526 => x"0c30c3",
   36527 => x"0c30c3",
   36528 => x"0c30c3",
   36529 => x"0c30c3",
   36530 => x"0c30c3",
   36531 => x"0c30c3",
   36532 => x"0c30c3",
   36533 => x"0c30c3",
   36534 => x"0c30c3",
   36535 => x"0c3aff",
   36536 => x"ffffff",
   36537 => x"ffffff",
   36538 => x"ffffff",
   36539 => x"ffffff",
   36540 => x"ffffff",
   36541 => x"ffffff",
   36542 => x"ffffff",
   36543 => x"ffffff",
   36544 => x"ffffff",
   36545 => x"ffffff",
   36546 => x"ffffff",
   36547 => x"ffffff",
   36548 => x"ffffff",
   36549 => x"fffa95",
   36550 => x"abffff",
   36551 => x"ffffff",
   36552 => x"ffffff",
   36553 => x"ffffff",
   36554 => x"ffffff",
   36555 => x"ffffff",
   36556 => x"ffffff",
   36557 => x"ffffff",
   36558 => x"ffffff",
   36559 => x"ffffff",
   36560 => x"ffffff",
   36561 => x"fffb8c",
   36562 => x"30c30c",
   36563 => x"30c30c",
   36564 => x"30c30c",
   36565 => x"30c30c",
   36566 => x"30c30c",
   36567 => x"30c30c",
   36568 => x"30c30c",
   36569 => x"30c30c",
   36570 => x"30c30c",
   36571 => x"30c30c",
   36572 => x"30c30c",
   36573 => x"208208",
   36574 => x"208208",
   36575 => x"208208",
   36576 => x"208208",
   36577 => x"208208",
   36578 => x"208208",
   36579 => x"208208",
   36580 => x"208208",
   36581 => x"208208",
   36582 => x"208208",
   36583 => x"208208",
   36584 => x"208208",
   36585 => x"208208",
   36586 => x"208208",
   36587 => x"208208",
   36588 => x"208208",
   36589 => x"208208",
   36590 => x"208208",
   36591 => x"208208",
   36592 => x"208208",
   36593 => x"208208",
   36594 => x"208208",
   36595 => x"208104",
   36596 => x"104104",
   36597 => x"104104",
   36598 => x"104104",
   36599 => x"104104",
   36600 => x"104104",
   36601 => x"104104",
   36602 => x"104104",
   36603 => x"104104",
   36604 => x"104104",
   36605 => x"104104",
   36606 => x"104104",
   36607 => x"104104",
   36608 => x"104104",
   36609 => x"104104",
   36610 => x"104104",
   36611 => x"104104",
   36612 => x"104104",
   36613 => x"104104",
   36614 => x"104104",
   36615 => x"104104",
   36616 => x"104104",
   36617 => x"104104",
   36618 => x"104000",
   36619 => x"000000",
   36620 => x"000000",
   36621 => x"000000",
   36622 => x"000000",
   36623 => x"000000",
   36624 => x"000000",
   36625 => x"000000",
   36626 => x"000000",
   36627 => x"000000",
   36628 => x"000000",
   36629 => x"00057f",
   36630 => x"ffffff",
   36631 => x"ffffff",
   36632 => x"ffffff",
   36633 => x"ffffff",
   36634 => x"ffffff",
   36635 => x"ffffff",
   36636 => x"ffffff",
   36637 => x"ffffff",
   36638 => x"ffffff",
   36639 => x"ffffff",
   36640 => x"ffffff",
   36641 => x"ffffff",
   36642 => x"ffffff",
   36643 => x"ffffff",
   36644 => x"ffffff",
   36645 => x"ffffff",
   36646 => x"ffffff",
   36647 => x"ffffff",
   36648 => x"ffffff",
   36649 => x"ffffff",
   36650 => x"ffffff",
   36651 => x"ffffff",
   36652 => x"ffffff",
   36653 => x"ac30c3",
   36654 => x"0c30c3",
   36655 => x"0c30c3",
   36656 => x"0c30c3",
   36657 => x"0c30c3",
   36658 => x"0c30c3",
   36659 => x"0c30c3",
   36660 => x"0c30c3",
   36661 => x"0c30c3",
   36662 => x"0c30c3",
   36663 => x"0c30c3",
   36664 => x"0c30c3",
   36665 => x"0c30c3",
   36666 => x"0c30c3",
   36667 => x"0c30c3",
   36668 => x"0c30c3",
   36669 => x"0c30c3",
   36670 => x"0c30c3",
   36671 => x"0c30c3",
   36672 => x"0c30c3",
   36673 => x"0c30c3",
   36674 => x"0c30c3",
   36675 => x"0c30c3",
   36676 => x"0c30c3",
   36677 => x"0c30c3",
   36678 => x"0c30c3",
   36679 => x"0c30c3",
   36680 => x"0c30c3",
   36681 => x"0c30c3",
   36682 => x"0c30c3",
   36683 => x"0c30c3",
   36684 => x"0c30c3",
   36685 => x"0c30c3",
   36686 => x"0c30c3",
   36687 => x"0c30c3",
   36688 => x"0c30c3",
   36689 => x"0c30c3",
   36690 => x"0c30c3",
   36691 => x"0c30c3",
   36692 => x"0c30c3",
   36693 => x"0c30c3",
   36694 => x"0c30c3",
   36695 => x"0d7fff",
   36696 => x"ffffff",
   36697 => x"ffffff",
   36698 => x"ffffff",
   36699 => x"ffffff",
   36700 => x"ffffff",
   36701 => x"ffffff",
   36702 => x"ffffff",
   36703 => x"ffffff",
   36704 => x"ffffff",
   36705 => x"ffffff",
   36706 => x"ffffff",
   36707 => x"ffffff",
   36708 => x"ffffff",
   36709 => x"fffa95",
   36710 => x"abffff",
   36711 => x"ffffff",
   36712 => x"ffffff",
   36713 => x"ffffff",
   36714 => x"ffffff",
   36715 => x"ffffff",
   36716 => x"ffffff",
   36717 => x"ffffff",
   36718 => x"ffffff",
   36719 => x"ffffff",
   36720 => x"ffffff",
   36721 => x"fffb8c",
   36722 => x"30c30c",
   36723 => x"30c30c",
   36724 => x"30c30c",
   36725 => x"30c30c",
   36726 => x"30c30c",
   36727 => x"30c30c",
   36728 => x"30c30c",
   36729 => x"30c30c",
   36730 => x"30c30c",
   36731 => x"30c30c",
   36732 => x"30c30c",
   36733 => x"208208",
   36734 => x"208208",
   36735 => x"208208",
   36736 => x"208208",
   36737 => x"208208",
   36738 => x"208208",
   36739 => x"208208",
   36740 => x"208208",
   36741 => x"208208",
   36742 => x"208208",
   36743 => x"208208",
   36744 => x"208208",
   36745 => x"208208",
   36746 => x"208208",
   36747 => x"208208",
   36748 => x"208208",
   36749 => x"208208",
   36750 => x"208208",
   36751 => x"208208",
   36752 => x"208208",
   36753 => x"208208",
   36754 => x"208208",
   36755 => x"208104",
   36756 => x"104104",
   36757 => x"104104",
   36758 => x"104104",
   36759 => x"104104",
   36760 => x"104104",
   36761 => x"104104",
   36762 => x"104104",
   36763 => x"104104",
   36764 => x"104104",
   36765 => x"104104",
   36766 => x"104104",
   36767 => x"104104",
   36768 => x"104104",
   36769 => x"104104",
   36770 => x"104104",
   36771 => x"104104",
   36772 => x"104104",
   36773 => x"104104",
   36774 => x"104104",
   36775 => x"104104",
   36776 => x"104104",
   36777 => x"104104",
   36778 => x"104000",
   36779 => x"000000",
   36780 => x"000000",
   36781 => x"000000",
   36782 => x"000000",
   36783 => x"000000",
   36784 => x"000000",
   36785 => x"000000",
   36786 => x"000000",
   36787 => x"000000",
   36788 => x"000000",
   36789 => x"00057f",
   36790 => x"ffffff",
   36791 => x"ffffff",
   36792 => x"ffffff",
   36793 => x"ffffff",
   36794 => x"ffffff",
   36795 => x"ffffff",
   36796 => x"ffffff",
   36797 => x"ffffff",
   36798 => x"ffffff",
   36799 => x"ffffff",
   36800 => x"ffffff",
   36801 => x"ffffff",
   36802 => x"ffffff",
   36803 => x"ffffff",
   36804 => x"ffffff",
   36805 => x"ffffff",
   36806 => x"ffffff",
   36807 => x"ffffff",
   36808 => x"ffffff",
   36809 => x"ffffff",
   36810 => x"ffffff",
   36811 => x"ffffff",
   36812 => x"ffffff",
   36813 => x"fd70c3",
   36814 => x"0c30c3",
   36815 => x"0c30c3",
   36816 => x"0c30c3",
   36817 => x"0c30c3",
   36818 => x"0c30c3",
   36819 => x"0c30c3",
   36820 => x"0c30c3",
   36821 => x"0c30c3",
   36822 => x"0c30c3",
   36823 => x"0c30c3",
   36824 => x"0c30c3",
   36825 => x"0c30c3",
   36826 => x"0c30c3",
   36827 => x"0c30c3",
   36828 => x"0c30c3",
   36829 => x"0c30c3",
   36830 => x"0c30c3",
   36831 => x"0c30c3",
   36832 => x"0c30c3",
   36833 => x"0c30c3",
   36834 => x"0c30c3",
   36835 => x"0c30c3",
   36836 => x"0c30c3",
   36837 => x"0c30c3",
   36838 => x"0c30c3",
   36839 => x"0c30c3",
   36840 => x"0c30c3",
   36841 => x"0c30c3",
   36842 => x"0c30c3",
   36843 => x"0c30c3",
   36844 => x"0c30c3",
   36845 => x"0c30c3",
   36846 => x"0c30c3",
   36847 => x"0c30c3",
   36848 => x"0c30c3",
   36849 => x"0c30c3",
   36850 => x"0c30c3",
   36851 => x"0c30c3",
   36852 => x"0c30c3",
   36853 => x"0c30c3",
   36854 => x"0c30c3",
   36855 => x"0ebfff",
   36856 => x"ffffff",
   36857 => x"ffffff",
   36858 => x"ffffff",
   36859 => x"ffffff",
   36860 => x"ffffff",
   36861 => x"ffffff",
   36862 => x"ffffff",
   36863 => x"ffffff",
   36864 => x"ffffff",
   36865 => x"ffffff",
   36866 => x"ffffff",
   36867 => x"ffffff",
   36868 => x"ffffff",
   36869 => x"fffa95",
   36870 => x"abffff",
   36871 => x"ffffff",
   36872 => x"ffffff",
   36873 => x"ffffff",
   36874 => x"ffffff",
   36875 => x"ffffff",
   36876 => x"ffffff",
   36877 => x"ffffff",
   36878 => x"ffffff",
   36879 => x"ffffff",
   36880 => x"ffffff",
   36881 => x"fffb8c",
   36882 => x"30c30c",
   36883 => x"30c30c",
   36884 => x"30c30c",
   36885 => x"30c30c",
   36886 => x"30c30c",
   36887 => x"30c30c",
   36888 => x"30c30c",
   36889 => x"30c30c",
   36890 => x"30c30c",
   36891 => x"30c30c",
   36892 => x"30c30c",
   36893 => x"208208",
   36894 => x"208208",
   36895 => x"208208",
   36896 => x"208208",
   36897 => x"208208",
   36898 => x"208208",
   36899 => x"208208",
   36900 => x"208208",
   36901 => x"208208",
   36902 => x"208208",
   36903 => x"208208",
   36904 => x"208208",
   36905 => x"208208",
   36906 => x"208208",
   36907 => x"208208",
   36908 => x"208208",
   36909 => x"208208",
   36910 => x"208208",
   36911 => x"208208",
   36912 => x"208208",
   36913 => x"208208",
   36914 => x"208208",
   36915 => x"208104",
   36916 => x"104104",
   36917 => x"104104",
   36918 => x"104104",
   36919 => x"104104",
   36920 => x"104104",
   36921 => x"104104",
   36922 => x"104104",
   36923 => x"104104",
   36924 => x"104104",
   36925 => x"104104",
   36926 => x"104104",
   36927 => x"104104",
   36928 => x"104104",
   36929 => x"104104",
   36930 => x"104104",
   36931 => x"104104",
   36932 => x"104104",
   36933 => x"104104",
   36934 => x"104104",
   36935 => x"104104",
   36936 => x"104104",
   36937 => x"104104",
   36938 => x"104000",
   36939 => x"000000",
   36940 => x"000000",
   36941 => x"000000",
   36942 => x"000000",
   36943 => x"000000",
   36944 => x"000000",
   36945 => x"000000",
   36946 => x"000000",
   36947 => x"000000",
   36948 => x"000000",
   36949 => x"00057f",
   36950 => x"ffffff",
   36951 => x"ffffff",
   36952 => x"ffffff",
   36953 => x"ffffff",
   36954 => x"ffffff",
   36955 => x"ffffff",
   36956 => x"fffaaa",
   36957 => x"aaaabf",
   36958 => x"ffffff",
   36959 => x"ffffff",
   36960 => x"ffffff",
   36961 => x"ffffff",
   36962 => x"ffffff",
   36963 => x"ffffff",
   36964 => x"ffffff",
   36965 => x"ffffff",
   36966 => x"ffffff",
   36967 => x"ffffff",
   36968 => x"ffffff",
   36969 => x"ffffff",
   36970 => x"ffffff",
   36971 => x"ffffff",
   36972 => x"ffffff",
   36973 => x"feb0c3",
   36974 => x"0c30c3",
   36975 => x"0c30c3",
   36976 => x"0c30c3",
   36977 => x"0c30c3",
   36978 => x"0c30c3",
   36979 => x"0c30c3",
   36980 => x"0c30c3",
   36981 => x"0c30c3",
   36982 => x"0c30c3",
   36983 => x"0c30c3",
   36984 => x"0c30c3",
   36985 => x"0c30c3",
   36986 => x"0c30c3",
   36987 => x"0c30c3",
   36988 => x"0c30c3",
   36989 => x"0c30c3",
   36990 => x"0c30c3",
   36991 => x"0c30c3",
   36992 => x"0c30c3",
   36993 => x"0c30c3",
   36994 => x"0c30c3",
   36995 => x"0c30c3",
   36996 => x"0c30c3",
   36997 => x"0c30c3",
   36998 => x"0c30c3",
   36999 => x"0c30c3",
   37000 => x"0c30c3",
   37001 => x"0c30c3",
   37002 => x"0c30c3",
   37003 => x"0c30c3",
   37004 => x"0c30c3",
   37005 => x"0c30c3",
   37006 => x"0c30c3",
   37007 => x"0c30c3",
   37008 => x"0c30c3",
   37009 => x"0c30c3",
   37010 => x"0c30c3",
   37011 => x"0c30c3",
   37012 => x"0c30c3",
   37013 => x"0c30c3",
   37014 => x"0c30c3",
   37015 => x"5fffff",
   37016 => x"ffffff",
   37017 => x"ffffff",
   37018 => x"ffffff",
   37019 => x"ffffff",
   37020 => x"ffffff",
   37021 => x"ffffff",
   37022 => x"ffffff",
   37023 => x"ffffff",
   37024 => x"ffffff",
   37025 => x"ffffff",
   37026 => x"ffffff",
   37027 => x"ffffff",
   37028 => x"ffffff",
   37029 => x"fffa95",
   37030 => x"abffff",
   37031 => x"ffffff",
   37032 => x"ffffff",
   37033 => x"ffffff",
   37034 => x"ffffff",
   37035 => x"ffffff",
   37036 => x"ffffff",
   37037 => x"ffffff",
   37038 => x"ffffff",
   37039 => x"ffffff",
   37040 => x"ffffff",
   37041 => x"fffb8c",
   37042 => x"30c30c",
   37043 => x"30c30c",
   37044 => x"30c30c",
   37045 => x"30c30c",
   37046 => x"30c30c",
   37047 => x"30c30c",
   37048 => x"30c30c",
   37049 => x"30c30c",
   37050 => x"30c30c",
   37051 => x"30c30c",
   37052 => x"30c30c",
   37053 => x"208208",
   37054 => x"208208",
   37055 => x"208208",
   37056 => x"208208",
   37057 => x"208208",
   37058 => x"208208",
   37059 => x"208208",
   37060 => x"208208",
   37061 => x"208208",
   37062 => x"208208",
   37063 => x"208208",
   37064 => x"208208",
   37065 => x"208208",
   37066 => x"208208",
   37067 => x"208208",
   37068 => x"208208",
   37069 => x"208208",
   37070 => x"208208",
   37071 => x"208208",
   37072 => x"208208",
   37073 => x"208208",
   37074 => x"208208",
   37075 => x"208104",
   37076 => x"104104",
   37077 => x"104104",
   37078 => x"104104",
   37079 => x"104104",
   37080 => x"104104",
   37081 => x"104104",
   37082 => x"104104",
   37083 => x"104104",
   37084 => x"104104",
   37085 => x"104104",
   37086 => x"104104",
   37087 => x"104104",
   37088 => x"104104",
   37089 => x"104104",
   37090 => x"104104",
   37091 => x"104104",
   37092 => x"104104",
   37093 => x"104104",
   37094 => x"104104",
   37095 => x"104104",
   37096 => x"104104",
   37097 => x"104104",
   37098 => x"104000",
   37099 => x"000000",
   37100 => x"000000",
   37101 => x"000000",
   37102 => x"000000",
   37103 => x"000000",
   37104 => x"000000",
   37105 => x"000000",
   37106 => x"000000",
   37107 => x"000000",
   37108 => x"000000",
   37109 => x"00057f",
   37110 => x"ffffff",
   37111 => x"ffffff",
   37112 => x"ffffff",
   37113 => x"ffffff",
   37114 => x"ffffff",
   37115 => x"fffaaa",
   37116 => x"555540",
   37117 => x"000015",
   37118 => x"555abf",
   37119 => x"ffffff",
   37120 => x"ffffff",
   37121 => x"ffffff",
   37122 => x"ffffff",
   37123 => x"ffffff",
   37124 => x"ffffff",
   37125 => x"ffffff",
   37126 => x"ffffff",
   37127 => x"ffffff",
   37128 => x"ffffff",
   37129 => x"ffffff",
   37130 => x"ffffff",
   37131 => x"ffffff",
   37132 => x"ffffff",
   37133 => x"fff5c3",
   37134 => x"0c30c3",
   37135 => x"0c30c3",
   37136 => x"0c30c3",
   37137 => x"0c30c3",
   37138 => x"0c30c3",
   37139 => x"0c30c3",
   37140 => x"0c30c3",
   37141 => x"0c30c3",
   37142 => x"0c30c3",
   37143 => x"0c30c3",
   37144 => x"0c30c3",
   37145 => x"0c30c3",
   37146 => x"0c30c3",
   37147 => x"0c30c3",
   37148 => x"0c30c3",
   37149 => x"0c30c3",
   37150 => x"0c30c3",
   37151 => x"0c30c3",
   37152 => x"0c30c3",
   37153 => x"0c30c3",
   37154 => x"0c30c3",
   37155 => x"0c30c3",
   37156 => x"0c30c3",
   37157 => x"0c30c3",
   37158 => x"0c30c3",
   37159 => x"0c30c3",
   37160 => x"0c30c3",
   37161 => x"0c30c3",
   37162 => x"0c30c3",
   37163 => x"0c30c3",
   37164 => x"0c30c3",
   37165 => x"0c30c3",
   37166 => x"0c30c3",
   37167 => x"0c30c3",
   37168 => x"0c30c3",
   37169 => x"0c30c3",
   37170 => x"0c30c3",
   37171 => x"0c30c3",
   37172 => x"0c30c3",
   37173 => x"0c30c3",
   37174 => x"0c30c3",
   37175 => x"afffff",
   37176 => x"ffffff",
   37177 => x"ffffff",
   37178 => x"ffffff",
   37179 => x"ffffff",
   37180 => x"ffffff",
   37181 => x"ffffff",
   37182 => x"ffffff",
   37183 => x"ffffff",
   37184 => x"ffffff",
   37185 => x"ffffff",
   37186 => x"ffffff",
   37187 => x"ffffff",
   37188 => x"ffffff",
   37189 => x"fffa95",
   37190 => x"abffff",
   37191 => x"ffffff",
   37192 => x"ffffff",
   37193 => x"ffffff",
   37194 => x"ffffff",
   37195 => x"ffffff",
   37196 => x"ffffff",
   37197 => x"ffffff",
   37198 => x"ffffff",
   37199 => x"ffffff",
   37200 => x"ffffff",
   37201 => x"fffb8c",
   37202 => x"30c30c",
   37203 => x"30c30c",
   37204 => x"30c30c",
   37205 => x"30c30c",
   37206 => x"30c30c",
   37207 => x"30c30c",
   37208 => x"30c30c",
   37209 => x"30c30c",
   37210 => x"30c30c",
   37211 => x"30c30c",
   37212 => x"30c30c",
   37213 => x"208208",
   37214 => x"208208",
   37215 => x"208208",
   37216 => x"208208",
   37217 => x"208208",
   37218 => x"208208",
   37219 => x"208208",
   37220 => x"208208",
   37221 => x"208208",
   37222 => x"208208",
   37223 => x"208208",
   37224 => x"208208",
   37225 => x"208208",
   37226 => x"208208",
   37227 => x"208208",
   37228 => x"208208",
   37229 => x"208208",
   37230 => x"208208",
   37231 => x"208208",
   37232 => x"208208",
   37233 => x"208208",
   37234 => x"208208",
   37235 => x"208104",
   37236 => x"104104",
   37237 => x"104104",
   37238 => x"104104",
   37239 => x"104104",
   37240 => x"104104",
   37241 => x"104104",
   37242 => x"104104",
   37243 => x"104104",
   37244 => x"104104",
   37245 => x"104104",
   37246 => x"104104",
   37247 => x"104104",
   37248 => x"104104",
   37249 => x"104104",
   37250 => x"104104",
   37251 => x"104104",
   37252 => x"104104",
   37253 => x"104104",
   37254 => x"104104",
   37255 => x"104104",
   37256 => x"104104",
   37257 => x"104104",
   37258 => x"104000",
   37259 => x"000000",
   37260 => x"000000",
   37261 => x"000000",
   37262 => x"000000",
   37263 => x"000000",
   37264 => x"000000",
   37265 => x"000000",
   37266 => x"000000",
   37267 => x"000000",
   37268 => x"000000",
   37269 => x"00057f",
   37270 => x"ffffff",
   37271 => x"ffffff",
   37272 => x"ffffff",
   37273 => x"ffffff",
   37274 => x"ffffff",
   37275 => x"a95000",
   37276 => x"000000",
   37277 => x"000000",
   37278 => x"000000",
   37279 => x"56afff",
   37280 => x"ffffff",
   37281 => x"ffffff",
   37282 => x"ffffff",
   37283 => x"ffffff",
   37284 => x"ffffff",
   37285 => x"ffffff",
   37286 => x"ffffff",
   37287 => x"ffffff",
   37288 => x"ffffff",
   37289 => x"ffffff",
   37290 => x"ffffff",
   37291 => x"ffffff",
   37292 => x"ffffff",
   37293 => x"fffac3",
   37294 => x"0c30c3",
   37295 => x"0c30c3",
   37296 => x"0c30c3",
   37297 => x"0c30c3",
   37298 => x"0c30c3",
   37299 => x"0c30c3",
   37300 => x"0c30c3",
   37301 => x"0c30c3",
   37302 => x"0c30c3",
   37303 => x"0c30c3",
   37304 => x"0c30c3",
   37305 => x"0c30c3",
   37306 => x"0c30c3",
   37307 => x"0c30c3",
   37308 => x"0c30c3",
   37309 => x"0c30c3",
   37310 => x"0c30c3",
   37311 => x"0c30c3",
   37312 => x"0c30c3",
   37313 => x"0c30c3",
   37314 => x"0c30c3",
   37315 => x"0c30c3",
   37316 => x"0c30c3",
   37317 => x"0c30c3",
   37318 => x"0c30c3",
   37319 => x"0c30c3",
   37320 => x"0c30c3",
   37321 => x"0c30c3",
   37322 => x"0c30c3",
   37323 => x"0c30c3",
   37324 => x"0c30c3",
   37325 => x"0c30c3",
   37326 => x"0c30c3",
   37327 => x"0c30c3",
   37328 => x"0c30c3",
   37329 => x"0c30c3",
   37330 => x"0c30c3",
   37331 => x"0c30c3",
   37332 => x"0c30c3",
   37333 => x"0c30c3",
   37334 => x"0c30d7",
   37335 => x"ffffff",
   37336 => x"ffffff",
   37337 => x"ffffff",
   37338 => x"ffffff",
   37339 => x"ffffff",
   37340 => x"ffffff",
   37341 => x"ffffff",
   37342 => x"ffffff",
   37343 => x"ffffff",
   37344 => x"ffffff",
   37345 => x"ffffff",
   37346 => x"ffffff",
   37347 => x"ffffff",
   37348 => x"ffffff",
   37349 => x"fffa95",
   37350 => x"abffff",
   37351 => x"ffffff",
   37352 => x"ffffff",
   37353 => x"ffffff",
   37354 => x"ffffff",
   37355 => x"ffffff",
   37356 => x"ffffff",
   37357 => x"ffffff",
   37358 => x"ffffff",
   37359 => x"ffffff",
   37360 => x"ffffff",
   37361 => x"fffb8c",
   37362 => x"30c30c",
   37363 => x"30c30c",
   37364 => x"30c30c",
   37365 => x"30c30c",
   37366 => x"30c30c",
   37367 => x"30c30c",
   37368 => x"30c30c",
   37369 => x"30c30c",
   37370 => x"30c30c",
   37371 => x"30c30c",
   37372 => x"30c30c",
   37373 => x"208208",
   37374 => x"208208",
   37375 => x"208208",
   37376 => x"208208",
   37377 => x"208208",
   37378 => x"208208",
   37379 => x"208208",
   37380 => x"208208",
   37381 => x"208208",
   37382 => x"208208",
   37383 => x"208208",
   37384 => x"208208",
   37385 => x"208208",
   37386 => x"208208",
   37387 => x"208208",
   37388 => x"208208",
   37389 => x"208208",
   37390 => x"208208",
   37391 => x"208208",
   37392 => x"208208",
   37393 => x"208208",
   37394 => x"208208",
   37395 => x"208104",
   37396 => x"104104",
   37397 => x"104104",
   37398 => x"104104",
   37399 => x"104104",
   37400 => x"104104",
   37401 => x"104104",
   37402 => x"104104",
   37403 => x"104104",
   37404 => x"104104",
   37405 => x"104104",
   37406 => x"104104",
   37407 => x"104104",
   37408 => x"104104",
   37409 => x"104104",
   37410 => x"104104",
   37411 => x"104104",
   37412 => x"104104",
   37413 => x"104104",
   37414 => x"104104",
   37415 => x"104104",
   37416 => x"104104",
   37417 => x"104104",
   37418 => x"104000",
   37419 => x"000000",
   37420 => x"000000",
   37421 => x"000000",
   37422 => x"000000",
   37423 => x"000000",
   37424 => x"000000",
   37425 => x"000000",
   37426 => x"000000",
   37427 => x"000000",
   37428 => x"000000",
   37429 => x"00057f",
   37430 => x"ffffff",
   37431 => x"ffffff",
   37432 => x"ffffff",
   37433 => x"ffffff",
   37434 => x"ffffd5",
   37435 => x"000000",
   37436 => x"000000",
   37437 => x"000000",
   37438 => x"000000",
   37439 => x"00057f",
   37440 => x"ffffff",
   37441 => x"ffffff",
   37442 => x"ffffff",
   37443 => x"ffffff",
   37444 => x"ffffff",
   37445 => x"ffffff",
   37446 => x"ffffff",
   37447 => x"ffffff",
   37448 => x"ffffff",
   37449 => x"ffffff",
   37450 => x"ffffff",
   37451 => x"ffffff",
   37452 => x"ffffff",
   37453 => x"ffffd7",
   37454 => x"0c30c3",
   37455 => x"0c30c3",
   37456 => x"0c30c3",
   37457 => x"0c30c3",
   37458 => x"0c30c3",
   37459 => x"0c30c3",
   37460 => x"0c30c3",
   37461 => x"0c30c3",
   37462 => x"0c30c3",
   37463 => x"0c30c3",
   37464 => x"0c30c3",
   37465 => x"0c30c3",
   37466 => x"0c30c3",
   37467 => x"0c30c3",
   37468 => x"0c30c3",
   37469 => x"0c30c3",
   37470 => x"0c30c3",
   37471 => x"0c30c3",
   37472 => x"0c30c3",
   37473 => x"0c30c3",
   37474 => x"0c30c3",
   37475 => x"0c30c3",
   37476 => x"0c30c3",
   37477 => x"0c30c3",
   37478 => x"0c30c3",
   37479 => x"0c30c3",
   37480 => x"0c30c3",
   37481 => x"0c30c3",
   37482 => x"0c30c3",
   37483 => x"0c30c3",
   37484 => x"0c30c3",
   37485 => x"0c30c3",
   37486 => x"0c30c3",
   37487 => x"0c30c3",
   37488 => x"0c30c3",
   37489 => x"0c30c3",
   37490 => x"0c30c3",
   37491 => x"0c30c3",
   37492 => x"0c30c3",
   37493 => x"0c30c3",
   37494 => x"0c30eb",
   37495 => x"ffffff",
   37496 => x"ffffff",
   37497 => x"ffffff",
   37498 => x"ffffff",
   37499 => x"ffffff",
   37500 => x"ffffff",
   37501 => x"ffffff",
   37502 => x"ffffff",
   37503 => x"ffffff",
   37504 => x"ffffff",
   37505 => x"ffffff",
   37506 => x"ffffff",
   37507 => x"ffffff",
   37508 => x"ffffff",
   37509 => x"fffa95",
   37510 => x"abffff",
   37511 => x"ffffff",
   37512 => x"ffffff",
   37513 => x"ffffff",
   37514 => x"ffffff",
   37515 => x"ffffff",
   37516 => x"ffffff",
   37517 => x"ffffff",
   37518 => x"ffffff",
   37519 => x"ffffff",
   37520 => x"ffffff",
   37521 => x"fffb8c",
   37522 => x"30c30c",
   37523 => x"30c30c",
   37524 => x"30c30c",
   37525 => x"30c30c",
   37526 => x"30c30c",
   37527 => x"30c30c",
   37528 => x"30c30c",
   37529 => x"30c30c",
   37530 => x"30c30c",
   37531 => x"30c30c",
   37532 => x"30c30c",
   37533 => x"208208",
   37534 => x"208208",
   37535 => x"208208",
   37536 => x"208208",
   37537 => x"208208",
   37538 => x"208208",
   37539 => x"208208",
   37540 => x"208208",
   37541 => x"208208",
   37542 => x"208208",
   37543 => x"208208",
   37544 => x"208208",
   37545 => x"208208",
   37546 => x"208208",
   37547 => x"208208",
   37548 => x"208208",
   37549 => x"208208",
   37550 => x"208208",
   37551 => x"208208",
   37552 => x"208208",
   37553 => x"208208",
   37554 => x"208208",
   37555 => x"208104",
   37556 => x"104104",
   37557 => x"104104",
   37558 => x"104104",
   37559 => x"104104",
   37560 => x"104104",
   37561 => x"104104",
   37562 => x"104104",
   37563 => x"104104",
   37564 => x"104104",
   37565 => x"104104",
   37566 => x"104104",
   37567 => x"104104",
   37568 => x"104104",
   37569 => x"104104",
   37570 => x"104104",
   37571 => x"104104",
   37572 => x"104104",
   37573 => x"104104",
   37574 => x"104104",
   37575 => x"104104",
   37576 => x"104104",
   37577 => x"104104",
   37578 => x"104000",
   37579 => x"000000",
   37580 => x"000000",
   37581 => x"000000",
   37582 => x"000000",
   37583 => x"000000",
   37584 => x"000000",
   37585 => x"000000",
   37586 => x"000000",
   37587 => x"000000",
   37588 => x"000000",
   37589 => x"00057f",
   37590 => x"ffffff",
   37591 => x"ffffff",
   37592 => x"ffffff",
   37593 => x"ffffff",
   37594 => x"fea540",
   37595 => x"000000",
   37596 => x"555aaa",
   37597 => x"aaaaaa",
   37598 => x"540000",
   37599 => x"00002a",
   37600 => x"ffffff",
   37601 => x"ffffff",
   37602 => x"ffffff",
   37603 => x"ffffff",
   37604 => x"ffffff",
   37605 => x"ffffff",
   37606 => x"ffffff",
   37607 => x"ffffff",
   37608 => x"ffffff",
   37609 => x"ffffff",
   37610 => x"ffffff",
   37611 => x"ffffff",
   37612 => x"ffffff",
   37613 => x"ffffeb",
   37614 => x"0c30c3",
   37615 => x"0c30c3",
   37616 => x"0c30c3",
   37617 => x"0c30c3",
   37618 => x"0c30c3",
   37619 => x"0c30c3",
   37620 => x"0c30c3",
   37621 => x"0c30c3",
   37622 => x"0c30c3",
   37623 => x"0c30c3",
   37624 => x"0c30c3",
   37625 => x"0c30c3",
   37626 => x"0c30c3",
   37627 => x"0c30c3",
   37628 => x"0c30c3",
   37629 => x"0c30c3",
   37630 => x"0c30c3",
   37631 => x"0c30c3",
   37632 => x"0c30c3",
   37633 => x"0c30c3",
   37634 => x"0c30c3",
   37635 => x"0c30c3",
   37636 => x"0c30c3",
   37637 => x"0c30c3",
   37638 => x"0c30c3",
   37639 => x"0c30c3",
   37640 => x"0c30c3",
   37641 => x"0c30c3",
   37642 => x"0c30c3",
   37643 => x"0c30c3",
   37644 => x"0c30c3",
   37645 => x"0c30c3",
   37646 => x"0c30c3",
   37647 => x"0c30c3",
   37648 => x"0c30c3",
   37649 => x"0c30c3",
   37650 => x"0c30c3",
   37651 => x"0c30c3",
   37652 => x"0c30c3",
   37653 => x"0c30c3",
   37654 => x"0c35ff",
   37655 => x"ffffff",
   37656 => x"ffffff",
   37657 => x"ffffff",
   37658 => x"ffffff",
   37659 => x"ffffff",
   37660 => x"ffffff",
   37661 => x"ffffff",
   37662 => x"ffffff",
   37663 => x"ffffff",
   37664 => x"ffffff",
   37665 => x"ffffff",
   37666 => x"ffffff",
   37667 => x"ffffff",
   37668 => x"ffffff",
   37669 => x"fffa95",
   37670 => x"abffff",
   37671 => x"ffffff",
   37672 => x"ffffff",
   37673 => x"ffffff",
   37674 => x"ffffff",
   37675 => x"ffffff",
   37676 => x"ffffff",
   37677 => x"ffffff",
   37678 => x"ffffff",
   37679 => x"ffffff",
   37680 => x"ffffff",
   37681 => x"fffb8c",
   37682 => x"30c30c",
   37683 => x"30c30c",
   37684 => x"30c30c",
   37685 => x"30c30c",
   37686 => x"30c30c",
   37687 => x"30c30c",
   37688 => x"30c30c",
   37689 => x"30c30c",
   37690 => x"30c30c",
   37691 => x"30c30c",
   37692 => x"30c30c",
   37693 => x"208208",
   37694 => x"208208",
   37695 => x"208208",
   37696 => x"208208",
   37697 => x"208208",
   37698 => x"208208",
   37699 => x"208208",
   37700 => x"208208",
   37701 => x"208208",
   37702 => x"208208",
   37703 => x"208208",
   37704 => x"208208",
   37705 => x"208208",
   37706 => x"208208",
   37707 => x"208208",
   37708 => x"208208",
   37709 => x"208208",
   37710 => x"208208",
   37711 => x"208208",
   37712 => x"208208",
   37713 => x"208208",
   37714 => x"208208",
   37715 => x"208104",
   37716 => x"104104",
   37717 => x"104104",
   37718 => x"104104",
   37719 => x"104104",
   37720 => x"104104",
   37721 => x"104104",
   37722 => x"104104",
   37723 => x"104104",
   37724 => x"104104",
   37725 => x"104104",
   37726 => x"104104",
   37727 => x"104104",
   37728 => x"104104",
   37729 => x"104104",
   37730 => x"104104",
   37731 => x"104104",
   37732 => x"104104",
   37733 => x"104104",
   37734 => x"104104",
   37735 => x"104104",
   37736 => x"104104",
   37737 => x"104104",
   37738 => x"104000",
   37739 => x"000000",
   37740 => x"000000",
   37741 => x"000000",
   37742 => x"000000",
   37743 => x"000000",
   37744 => x"000000",
   37745 => x"000000",
   37746 => x"000000",
   37747 => x"000000",
   37748 => x"000000",
   37749 => x"00057f",
   37750 => x"ffffff",
   37751 => x"ffffff",
   37752 => x"ffffff",
   37753 => x"ffffff",
   37754 => x"fd5000",
   37755 => x"00056a",
   37756 => x"ffffff",
   37757 => x"ffffff",
   37758 => x"fffa95",
   37759 => x"00002a",
   37760 => x"ffffff",
   37761 => x"ffffff",
   37762 => x"ffffff",
   37763 => x"ffffff",
   37764 => x"ffffff",
   37765 => x"ffffff",
   37766 => x"ffffff",
   37767 => x"ffffff",
   37768 => x"ffffff",
   37769 => x"ffffff",
   37770 => x"ffffff",
   37771 => x"ffffff",
   37772 => x"ffffff",
   37773 => x"ffffff",
   37774 => x"5c30c3",
   37775 => x"0c30c3",
   37776 => x"0c30c3",
   37777 => x"0c30c3",
   37778 => x"0c30c3",
   37779 => x"0c30c3",
   37780 => x"0c30c3",
   37781 => x"0c30c3",
   37782 => x"0c30c3",
   37783 => x"0c30c3",
   37784 => x"0c30c3",
   37785 => x"0c30c3",
   37786 => x"0c30c3",
   37787 => x"0c30c3",
   37788 => x"0c30c3",
   37789 => x"0c30c3",
   37790 => x"0c30c3",
   37791 => x"0c30c3",
   37792 => x"0c30c3",
   37793 => x"0c30c3",
   37794 => x"0c30c3",
   37795 => x"0c30c3",
   37796 => x"0c30c3",
   37797 => x"0c30c3",
   37798 => x"0c30c3",
   37799 => x"0c30c3",
   37800 => x"0c30c3",
   37801 => x"0c30c3",
   37802 => x"0c30c3",
   37803 => x"0c30c3",
   37804 => x"0c30c3",
   37805 => x"0c30c3",
   37806 => x"0c30c3",
   37807 => x"0c30c3",
   37808 => x"0c30c3",
   37809 => x"0c30c3",
   37810 => x"0c30c3",
   37811 => x"0c30c3",
   37812 => x"0c30c3",
   37813 => x"0c30c3",
   37814 => x"0c3aff",
   37815 => x"ffffff",
   37816 => x"ffffff",
   37817 => x"ffffff",
   37818 => x"ffffff",
   37819 => x"ffffff",
   37820 => x"ffffff",
   37821 => x"ffffff",
   37822 => x"ffffff",
   37823 => x"ffffff",
   37824 => x"ffffff",
   37825 => x"ffffff",
   37826 => x"ffffff",
   37827 => x"ffffff",
   37828 => x"ffffff",
   37829 => x"fffa95",
   37830 => x"abffff",
   37831 => x"ffffff",
   37832 => x"ffffff",
   37833 => x"ffffff",
   37834 => x"ffffff",
   37835 => x"ffffff",
   37836 => x"ffffff",
   37837 => x"ffffff",
   37838 => x"ffffff",
   37839 => x"ffffff",
   37840 => x"ffffff",
   37841 => x"fffb8c",
   37842 => x"30c30c",
   37843 => x"30c30c",
   37844 => x"30c30c",
   37845 => x"30c30c",
   37846 => x"30c30c",
   37847 => x"30c30c",
   37848 => x"30c30c",
   37849 => x"30c30c",
   37850 => x"30c30c",
   37851 => x"30c30c",
   37852 => x"30c30c",
   37853 => x"208208",
   37854 => x"208208",
   37855 => x"208208",
   37856 => x"208208",
   37857 => x"208208",
   37858 => x"208208",
   37859 => x"208208",
   37860 => x"208208",
   37861 => x"208208",
   37862 => x"208208",
   37863 => x"208208",
   37864 => x"208208",
   37865 => x"208208",
   37866 => x"208208",
   37867 => x"208208",
   37868 => x"208208",
   37869 => x"208208",
   37870 => x"208208",
   37871 => x"208208",
   37872 => x"208208",
   37873 => x"208208",
   37874 => x"208208",
   37875 => x"208104",
   37876 => x"104104",
   37877 => x"104104",
   37878 => x"104104",
   37879 => x"104104",
   37880 => x"104104",
   37881 => x"104104",
   37882 => x"104104",
   37883 => x"104104",
   37884 => x"104104",
   37885 => x"104104",
   37886 => x"104104",
   37887 => x"104104",
   37888 => x"104104",
   37889 => x"104104",
   37890 => x"104104",
   37891 => x"104104",
   37892 => x"104104",
   37893 => x"104104",
   37894 => x"104104",
   37895 => x"104104",
   37896 => x"104104",
   37897 => x"104104",
   37898 => x"104000",
   37899 => x"000000",
   37900 => x"000000",
   37901 => x"000000",
   37902 => x"000000",
   37903 => x"000000",
   37904 => x"000000",
   37905 => x"000000",
   37906 => x"000000",
   37907 => x"000000",
   37908 => x"000000",
   37909 => x"00057f",
   37910 => x"ffffff",
   37911 => x"ffffff",
   37912 => x"ffffff",
   37913 => x"ffffff",
   37914 => x"540000",
   37915 => x"015fff",
   37916 => x"ffffff",
   37917 => x"ffffff",
   37918 => x"ffffff",
   37919 => x"a9502a",
   37920 => x"ffffff",
   37921 => x"ffffff",
   37922 => x"ffffff",
   37923 => x"ffffff",
   37924 => x"ffffff",
   37925 => x"ffffff",
   37926 => x"ffffff",
   37927 => x"ffffff",
   37928 => x"ffffff",
   37929 => x"ffffff",
   37930 => x"ffffff",
   37931 => x"ffffff",
   37932 => x"ffffff",
   37933 => x"ffffff",
   37934 => x"ac30c3",
   37935 => x"0c30c3",
   37936 => x"0c30c3",
   37937 => x"0c30c3",
   37938 => x"0c30c3",
   37939 => x"0c30c3",
   37940 => x"0c30c3",
   37941 => x"0c30c3",
   37942 => x"0c30c3",
   37943 => x"0c30c3",
   37944 => x"0c30c3",
   37945 => x"0c30c3",
   37946 => x"0c30c3",
   37947 => x"0c30c3",
   37948 => x"0c30c3",
   37949 => x"0c30c3",
   37950 => x"0c30c3",
   37951 => x"0c30c3",
   37952 => x"0c30c3",
   37953 => x"0c30c3",
   37954 => x"0c30c3",
   37955 => x"0c30c3",
   37956 => x"0c30c3",
   37957 => x"0c30c3",
   37958 => x"0c30c3",
   37959 => x"0c30c3",
   37960 => x"0c30c3",
   37961 => x"0c30c3",
   37962 => x"0c30c3",
   37963 => x"0c30c3",
   37964 => x"0c30c3",
   37965 => x"0c30c3",
   37966 => x"0c30c3",
   37967 => x"0c30c3",
   37968 => x"0c30c3",
   37969 => x"0c30c3",
   37970 => x"0c30c3",
   37971 => x"0c30c3",
   37972 => x"0c30c3",
   37973 => x"0c30c3",
   37974 => x"0d7fff",
   37975 => x"ffffff",
   37976 => x"ffffff",
   37977 => x"ffffff",
   37978 => x"ffffff",
   37979 => x"ffffff",
   37980 => x"ffffff",
   37981 => x"ffffff",
   37982 => x"ffffff",
   37983 => x"ffffff",
   37984 => x"ffffff",
   37985 => x"ffffff",
   37986 => x"ffffff",
   37987 => x"ffffff",
   37988 => x"ffffff",
   37989 => x"fffa95",
   37990 => x"abffff",
   37991 => x"ffffff",
   37992 => x"ffffff",
   37993 => x"ffffff",
   37994 => x"ffffff",
   37995 => x"ffffff",
   37996 => x"ffffff",
   37997 => x"ffffff",
   37998 => x"ffffff",
   37999 => x"ffffff",
   38000 => x"ffffff",
   38001 => x"fffb8c",
   38002 => x"30c30c",
   38003 => x"30c30c",
   38004 => x"30c30c",
   38005 => x"30c30c",
   38006 => x"30c30c",
   38007 => x"30c30c",
   38008 => x"30c30c",
   38009 => x"30c30c",
   38010 => x"30c30c",
   38011 => x"30c30c",
   38012 => x"30c30c",
   38013 => x"208208",
   38014 => x"208208",
   38015 => x"208208",
   38016 => x"208208",
   38017 => x"208208",
   38018 => x"208208",
   38019 => x"208208",
   38020 => x"208208",
   38021 => x"208208",
   38022 => x"208208",
   38023 => x"208208",
   38024 => x"208208",
   38025 => x"208208",
   38026 => x"208208",
   38027 => x"208208",
   38028 => x"208208",
   38029 => x"208208",
   38030 => x"208208",
   38031 => x"208208",
   38032 => x"208208",
   38033 => x"208208",
   38034 => x"208208",
   38035 => x"208104",
   38036 => x"104104",
   38037 => x"104104",
   38038 => x"104104",
   38039 => x"104104",
   38040 => x"104104",
   38041 => x"104104",
   38042 => x"104104",
   38043 => x"104104",
   38044 => x"104104",
   38045 => x"104104",
   38046 => x"104104",
   38047 => x"104104",
   38048 => x"104104",
   38049 => x"104104",
   38050 => x"104104",
   38051 => x"104104",
   38052 => x"104104",
   38053 => x"104104",
   38054 => x"104104",
   38055 => x"104104",
   38056 => x"104104",
   38057 => x"104104",
   38058 => x"104000",
   38059 => x"000000",
   38060 => x"000000",
   38061 => x"000000",
   38062 => x"000000",
   38063 => x"000000",
   38064 => x"000000",
   38065 => x"000000",
   38066 => x"000000",
   38067 => x"000000",
   38068 => x"000000",
   38069 => x"00057f",
   38070 => x"ffffff",
   38071 => x"ffffff",
   38072 => x"ffffff",
   38073 => x"ffffea",
   38074 => x"000000",
   38075 => x"abffff",
   38076 => x"ffffff",
   38077 => x"ffffff",
   38078 => x"ffffff",
   38079 => x"fffaaa",
   38080 => x"ffffff",
   38081 => x"ffffff",
   38082 => x"ffffff",
   38083 => x"ffffff",
   38084 => x"ffffff",
   38085 => x"ffffff",
   38086 => x"ffffff",
   38087 => x"ffffff",
   38088 => x"ffffff",
   38089 => x"ffffff",
   38090 => x"ffffff",
   38091 => x"ffffff",
   38092 => x"ffffff",
   38093 => x"ffffff",
   38094 => x"feb0c3",
   38095 => x"0c30c3",
   38096 => x"0c30c3",
   38097 => x"0c30c3",
   38098 => x"0c30c3",
   38099 => x"0c30c3",
   38100 => x"0c30c3",
   38101 => x"0c30c3",
   38102 => x"0c30c3",
   38103 => x"0c30c3",
   38104 => x"0c30c3",
   38105 => x"0c30c3",
   38106 => x"0c30c3",
   38107 => x"0c30c3",
   38108 => x"0c30c3",
   38109 => x"0c30c3",
   38110 => x"0c30c3",
   38111 => x"0c30c3",
   38112 => x"0c30c3",
   38113 => x"0c30c3",
   38114 => x"0c30c3",
   38115 => x"0c30c3",
   38116 => x"0c30c3",
   38117 => x"0c30c3",
   38118 => x"0c30c3",
   38119 => x"0c30c3",
   38120 => x"0c30c3",
   38121 => x"0c30c3",
   38122 => x"0c30c3",
   38123 => x"0c30c3",
   38124 => x"0c30c3",
   38125 => x"0c30c3",
   38126 => x"0c30c3",
   38127 => x"0c30c3",
   38128 => x"0c30c3",
   38129 => x"0c30c3",
   38130 => x"0c30c3",
   38131 => x"0c30c3",
   38132 => x"0c30c3",
   38133 => x"0c30c3",
   38134 => x"0ebfff",
   38135 => x"ffffff",
   38136 => x"ffffff",
   38137 => x"ffffff",
   38138 => x"ffffff",
   38139 => x"ffffff",
   38140 => x"ffffff",
   38141 => x"ffffff",
   38142 => x"ffffff",
   38143 => x"ffffff",
   38144 => x"ffffff",
   38145 => x"ffffff",
   38146 => x"ffffff",
   38147 => x"ffffff",
   38148 => x"ffffff",
   38149 => x"fffa95",
   38150 => x"abffff",
   38151 => x"ffffff",
   38152 => x"ffffff",
   38153 => x"ffffff",
   38154 => x"ffffff",
   38155 => x"ffffff",
   38156 => x"ffffff",
   38157 => x"ffffff",
   38158 => x"ffffff",
   38159 => x"ffffff",
   38160 => x"ffffff",
   38161 => x"fffb8c",
   38162 => x"30c30c",
   38163 => x"30c30c",
   38164 => x"30c30c",
   38165 => x"30c30c",
   38166 => x"30c30c",
   38167 => x"30c30c",
   38168 => x"30c30c",
   38169 => x"30c30c",
   38170 => x"30c30c",
   38171 => x"30c30c",
   38172 => x"30c30c",
   38173 => x"208208",
   38174 => x"208208",
   38175 => x"208208",
   38176 => x"208208",
   38177 => x"208208",
   38178 => x"208208",
   38179 => x"208208",
   38180 => x"208208",
   38181 => x"208208",
   38182 => x"208208",
   38183 => x"208208",
   38184 => x"208208",
   38185 => x"208208",
   38186 => x"208208",
   38187 => x"208208",
   38188 => x"208208",
   38189 => x"208208",
   38190 => x"208208",
   38191 => x"208208",
   38192 => x"208208",
   38193 => x"208208",
   38194 => x"208208",
   38195 => x"208104",
   38196 => x"104104",
   38197 => x"104104",
   38198 => x"104104",
   38199 => x"104104",
   38200 => x"104104",
   38201 => x"104104",
   38202 => x"104104",
   38203 => x"104104",
   38204 => x"104104",
   38205 => x"104104",
   38206 => x"104104",
   38207 => x"104104",
   38208 => x"104104",
   38209 => x"104104",
   38210 => x"104104",
   38211 => x"104104",
   38212 => x"104104",
   38213 => x"104104",
   38214 => x"104104",
   38215 => x"104104",
   38216 => x"104104",
   38217 => x"104104",
   38218 => x"104000",
   38219 => x"000000",
   38220 => x"000000",
   38221 => x"000000",
   38222 => x"000000",
   38223 => x"000000",
   38224 => x"000000",
   38225 => x"000000",
   38226 => x"000000",
   38227 => x"000000",
   38228 => x"000000",
   38229 => x"00057f",
   38230 => x"ffffff",
   38231 => x"ffffff",
   38232 => x"ffffff",
   38233 => x"ffffd5",
   38234 => x"000015",
   38235 => x"ffffff",
   38236 => x"ffffff",
   38237 => x"ffffff",
   38238 => x"ffffff",
   38239 => x"ffffff",
   38240 => x"ffffff",
   38241 => x"ffffff",
   38242 => x"ffffff",
   38243 => x"ffffff",
   38244 => x"ffffff",
   38245 => x"ffffff",
   38246 => x"ffffff",
   38247 => x"ffffff",
   38248 => x"ffffff",
   38249 => x"ffffff",
   38250 => x"ffffff",
   38251 => x"ffffff",
   38252 => x"ffffff",
   38253 => x"ffffff",
   38254 => x"fff5c3",
   38255 => x"0c30c3",
   38256 => x"0c30c3",
   38257 => x"0c30c3",
   38258 => x"0c30c3",
   38259 => x"0c30c3",
   38260 => x"0c30c3",
   38261 => x"0c30c3",
   38262 => x"0c30c3",
   38263 => x"0c30c3",
   38264 => x"0c30c3",
   38265 => x"0c30c3",
   38266 => x"0c30c3",
   38267 => x"0c30c3",
   38268 => x"0c30c3",
   38269 => x"0c30c3",
   38270 => x"0c30c3",
   38271 => x"0c30c3",
   38272 => x"0c30c3",
   38273 => x"0c30c3",
   38274 => x"0c30c3",
   38275 => x"0c30c3",
   38276 => x"0c30c3",
   38277 => x"0c30c3",
   38278 => x"0c30c3",
   38279 => x"0c30c3",
   38280 => x"0c30c3",
   38281 => x"0c30c3",
   38282 => x"0c30c3",
   38283 => x"0c30c3",
   38284 => x"0c30c3",
   38285 => x"0c30c3",
   38286 => x"0c30c3",
   38287 => x"0c30c3",
   38288 => x"0c30c3",
   38289 => x"0c30c3",
   38290 => x"0c30c3",
   38291 => x"0c30c3",
   38292 => x"0c30c3",
   38293 => x"0c30c3",
   38294 => x"afffff",
   38295 => x"ffffff",
   38296 => x"ffffff",
   38297 => x"ffffff",
   38298 => x"ffffff",
   38299 => x"ffffff",
   38300 => x"ffffff",
   38301 => x"ffffff",
   38302 => x"ffffff",
   38303 => x"ffffff",
   38304 => x"ffffff",
   38305 => x"ffffff",
   38306 => x"ffffff",
   38307 => x"ffffff",
   38308 => x"ffffff",
   38309 => x"fffa95",
   38310 => x"abffff",
   38311 => x"ffffff",
   38312 => x"ffffff",
   38313 => x"ffffff",
   38314 => x"ffffff",
   38315 => x"ffffff",
   38316 => x"ffffff",
   38317 => x"ffffff",
   38318 => x"ffffff",
   38319 => x"ffffff",
   38320 => x"ffffff",
   38321 => x"fffb8c",
   38322 => x"30c30c",
   38323 => x"30c30c",
   38324 => x"30c30c",
   38325 => x"30c30c",
   38326 => x"30c30c",
   38327 => x"30c30c",
   38328 => x"30c30c",
   38329 => x"30c30c",
   38330 => x"30c30c",
   38331 => x"30c30c",
   38332 => x"30c30c",
   38333 => x"208208",
   38334 => x"208208",
   38335 => x"208208",
   38336 => x"208208",
   38337 => x"208208",
   38338 => x"208208",
   38339 => x"208208",
   38340 => x"208208",
   38341 => x"208208",
   38342 => x"208208",
   38343 => x"208208",
   38344 => x"208208",
   38345 => x"208208",
   38346 => x"208208",
   38347 => x"208208",
   38348 => x"208208",
   38349 => x"208208",
   38350 => x"208208",
   38351 => x"208208",
   38352 => x"208208",
   38353 => x"208208",
   38354 => x"208208",
   38355 => x"208104",
   38356 => x"104104",
   38357 => x"104104",
   38358 => x"104104",
   38359 => x"104104",
   38360 => x"104104",
   38361 => x"104104",
   38362 => x"104104",
   38363 => x"104104",
   38364 => x"104104",
   38365 => x"104104",
   38366 => x"104104",
   38367 => x"104104",
   38368 => x"104104",
   38369 => x"104104",
   38370 => x"104104",
   38371 => x"104104",
   38372 => x"104104",
   38373 => x"104104",
   38374 => x"104104",
   38375 => x"104104",
   38376 => x"104104",
   38377 => x"104104",
   38378 => x"104000",
   38379 => x"000000",
   38380 => x"000000",
   38381 => x"000000",
   38382 => x"000000",
   38383 => x"000000",
   38384 => x"000000",
   38385 => x"000000",
   38386 => x"000000",
   38387 => x"000000",
   38388 => x"000000",
   38389 => x"00057f",
   38390 => x"ffffff",
   38391 => x"ffffff",
   38392 => x"ffffff",
   38393 => x"fffa80",
   38394 => x"00002a",
   38395 => x"ffffff",
   38396 => x"ffffff",
   38397 => x"ffffff",
   38398 => x"ffffff",
   38399 => x"ffffff",
   38400 => x"ffffff",
   38401 => x"ffffff",
   38402 => x"ffffff",
   38403 => x"ffffff",
   38404 => x"ffffff",
   38405 => x"ffffff",
   38406 => x"ffffff",
   38407 => x"ffffff",
   38408 => x"ffffff",
   38409 => x"ffffff",
   38410 => x"ffffff",
   38411 => x"ffffff",
   38412 => x"ffffff",
   38413 => x"ffffff",
   38414 => x"fffac3",
   38415 => x"0c30c3",
   38416 => x"0c30c3",
   38417 => x"0c30c3",
   38418 => x"0c30c3",
   38419 => x"0c30c3",
   38420 => x"0c30c3",
   38421 => x"0c30c3",
   38422 => x"0c30c3",
   38423 => x"0c30c3",
   38424 => x"0c30c3",
   38425 => x"0c30c3",
   38426 => x"0c30c3",
   38427 => x"0c30c3",
   38428 => x"0c30c3",
   38429 => x"0c30c3",
   38430 => x"0c30c3",
   38431 => x"0c30c3",
   38432 => x"0c30c3",
   38433 => x"0c30c3",
   38434 => x"0c30c3",
   38435 => x"0c30c3",
   38436 => x"0c30c3",
   38437 => x"0c30c3",
   38438 => x"0c30c3",
   38439 => x"0c30c3",
   38440 => x"0c30c3",
   38441 => x"0c30c3",
   38442 => x"0c30c3",
   38443 => x"0c30c3",
   38444 => x"0c30c3",
   38445 => x"0c30c3",
   38446 => x"0c30c3",
   38447 => x"0c30c3",
   38448 => x"0c30c3",
   38449 => x"0c30c3",
   38450 => x"0c30c3",
   38451 => x"0c30c3",
   38452 => x"0c30c3",
   38453 => x"0c30d7",
   38454 => x"ffffff",
   38455 => x"ffffff",
   38456 => x"ffffff",
   38457 => x"ffffff",
   38458 => x"ffffff",
   38459 => x"ffffff",
   38460 => x"ffffff",
   38461 => x"ffffff",
   38462 => x"ffffff",
   38463 => x"ffffff",
   38464 => x"ffffff",
   38465 => x"ffffff",
   38466 => x"ffffff",
   38467 => x"ffffff",
   38468 => x"ffffff",
   38469 => x"fffa95",
   38470 => x"abffff",
   38471 => x"ffffff",
   38472 => x"ffffff",
   38473 => x"ffffff",
   38474 => x"ffffff",
   38475 => x"ffffff",
   38476 => x"ffffff",
   38477 => x"ffffff",
   38478 => x"ffffff",
   38479 => x"ffffff",
   38480 => x"ffffff",
   38481 => x"fffb8c",
   38482 => x"30c30c",
   38483 => x"30c30c",
   38484 => x"30c30c",
   38485 => x"30c30c",
   38486 => x"30c30c",
   38487 => x"30c30c",
   38488 => x"30c30c",
   38489 => x"30c30c",
   38490 => x"30c30c",
   38491 => x"30c30c",
   38492 => x"30c30c",
   38493 => x"208208",
   38494 => x"208208",
   38495 => x"208208",
   38496 => x"208208",
   38497 => x"208208",
   38498 => x"208208",
   38499 => x"208208",
   38500 => x"208208",
   38501 => x"208208",
   38502 => x"208208",
   38503 => x"208208",
   38504 => x"208208",
   38505 => x"208208",
   38506 => x"208208",
   38507 => x"208208",
   38508 => x"208208",
   38509 => x"208208",
   38510 => x"208208",
   38511 => x"208208",
   38512 => x"208208",
   38513 => x"208208",
   38514 => x"208208",
   38515 => x"208104",
   38516 => x"104104",
   38517 => x"104104",
   38518 => x"104104",
   38519 => x"104104",
   38520 => x"104104",
   38521 => x"104104",
   38522 => x"104104",
   38523 => x"104104",
   38524 => x"104104",
   38525 => x"104104",
   38526 => x"104104",
   38527 => x"104104",
   38528 => x"104104",
   38529 => x"104104",
   38530 => x"104104",
   38531 => x"104104",
   38532 => x"104104",
   38533 => x"104104",
   38534 => x"104104",
   38535 => x"104104",
   38536 => x"104104",
   38537 => x"104104",
   38538 => x"104000",
   38539 => x"000000",
   38540 => x"000000",
   38541 => x"000000",
   38542 => x"000000",
   38543 => x"000000",
   38544 => x"000000",
   38545 => x"000000",
   38546 => x"000000",
   38547 => x"000000",
   38548 => x"000000",
   38549 => x"00057f",
   38550 => x"ffffff",
   38551 => x"ffffff",
   38552 => x"ffffff",
   38553 => x"fff540",
   38554 => x"00057f",
   38555 => x"ffffff",
   38556 => x"ffffff",
   38557 => x"ffffff",
   38558 => x"ffffff",
   38559 => x"ffffff",
   38560 => x"ffffff",
   38561 => x"ffffff",
   38562 => x"ffffff",
   38563 => x"ffffff",
   38564 => x"ffffff",
   38565 => x"ffffff",
   38566 => x"ffffff",
   38567 => x"ffffff",
   38568 => x"ffffff",
   38569 => x"ffffff",
   38570 => x"ffffff",
   38571 => x"ffffff",
   38572 => x"ffffff",
   38573 => x"ffffff",
   38574 => x"ffffd7",
   38575 => x"0c30c3",
   38576 => x"0c30c3",
   38577 => x"0c30c3",
   38578 => x"0c30c3",
   38579 => x"0c30c3",
   38580 => x"0c30c3",
   38581 => x"0c30c3",
   38582 => x"0c30c3",
   38583 => x"0c30c3",
   38584 => x"0c30c3",
   38585 => x"0c30c3",
   38586 => x"0c30c3",
   38587 => x"0c30c3",
   38588 => x"0c30c3",
   38589 => x"0c30c3",
   38590 => x"0c30c3",
   38591 => x"0c30c3",
   38592 => x"0c30c3",
   38593 => x"0c30c3",
   38594 => x"0c30c3",
   38595 => x"0c30c3",
   38596 => x"0c30c3",
   38597 => x"0c30c3",
   38598 => x"0c30c3",
   38599 => x"0c30c3",
   38600 => x"0c30c3",
   38601 => x"0c30c3",
   38602 => x"0c30c3",
   38603 => x"0c30c3",
   38604 => x"0c30c3",
   38605 => x"0c30c3",
   38606 => x"0c30c3",
   38607 => x"0c30c3",
   38608 => x"0c30c3",
   38609 => x"0c30c3",
   38610 => x"0c30c3",
   38611 => x"0c30c3",
   38612 => x"0c30c3",
   38613 => x"0c30eb",
   38614 => x"ffffff",
   38615 => x"ffffff",
   38616 => x"ffffff",
   38617 => x"ffffff",
   38618 => x"ffffff",
   38619 => x"ffffff",
   38620 => x"ffffff",
   38621 => x"ffffff",
   38622 => x"ffffff",
   38623 => x"ffffff",
   38624 => x"ffffff",
   38625 => x"ffffff",
   38626 => x"ffffff",
   38627 => x"ffffff",
   38628 => x"ffffff",
   38629 => x"fffa95",
   38630 => x"abffff",
   38631 => x"ffffff",
   38632 => x"ffffff",
   38633 => x"ffffff",
   38634 => x"ffffff",
   38635 => x"ffffff",
   38636 => x"ffffff",
   38637 => x"ffffff",
   38638 => x"ffffff",
   38639 => x"ffffff",
   38640 => x"ffffff",
   38641 => x"fffb8c",
   38642 => x"30c30c",
   38643 => x"30c30c",
   38644 => x"30c30c",
   38645 => x"30c30c",
   38646 => x"30c30c",
   38647 => x"30c30c",
   38648 => x"30c30c",
   38649 => x"30c30c",
   38650 => x"30c30c",
   38651 => x"30c30c",
   38652 => x"30c30c",
   38653 => x"208208",
   38654 => x"208208",
   38655 => x"208208",
   38656 => x"208208",
   38657 => x"208208",
   38658 => x"208208",
   38659 => x"208208",
   38660 => x"208208",
   38661 => x"208208",
   38662 => x"208208",
   38663 => x"208208",
   38664 => x"208208",
   38665 => x"208208",
   38666 => x"208208",
   38667 => x"208208",
   38668 => x"208208",
   38669 => x"208208",
   38670 => x"208208",
   38671 => x"208208",
   38672 => x"208208",
   38673 => x"208208",
   38674 => x"208208",
   38675 => x"208104",
   38676 => x"104104",
   38677 => x"104104",
   38678 => x"104104",
   38679 => x"104104",
   38680 => x"104104",
   38681 => x"104104",
   38682 => x"104104",
   38683 => x"104104",
   38684 => x"104104",
   38685 => x"104104",
   38686 => x"104104",
   38687 => x"104104",
   38688 => x"104104",
   38689 => x"104104",
   38690 => x"104104",
   38691 => x"104104",
   38692 => x"104104",
   38693 => x"104104",
   38694 => x"104104",
   38695 => x"104104",
   38696 => x"104104",
   38697 => x"104104",
   38698 => x"104000",
   38699 => x"000000",
   38700 => x"000000",
   38701 => x"000000",
   38702 => x"000000",
   38703 => x"000000",
   38704 => x"000000",
   38705 => x"000000",
   38706 => x"000000",
   38707 => x"000000",
   38708 => x"000000",
   38709 => x"00057f",
   38710 => x"ffffff",
   38711 => x"ffffff",
   38712 => x"ffffff",
   38713 => x"fff540",
   38714 => x"000abf",
   38715 => x"ffffff",
   38716 => x"ffffff",
   38717 => x"ffffff",
   38718 => x"ffffff",
   38719 => x"ffffff",
   38720 => x"ffffff",
   38721 => x"ffffff",
   38722 => x"ffffff",
   38723 => x"ffffff",
   38724 => x"ffffff",
   38725 => x"ffffff",
   38726 => x"ffffff",
   38727 => x"ffffff",
   38728 => x"ffffff",
   38729 => x"ffffff",
   38730 => x"ffffff",
   38731 => x"ffffff",
   38732 => x"ffffff",
   38733 => x"ffffff",
   38734 => x"ffffeb",
   38735 => x"5c30c3",
   38736 => x"0c30c3",
   38737 => x"0c30c3",
   38738 => x"0c30c3",
   38739 => x"0c30c3",
   38740 => x"0c30c3",
   38741 => x"0c30c3",
   38742 => x"0c30c3",
   38743 => x"0c30c3",
   38744 => x"0c30c3",
   38745 => x"0c30c3",
   38746 => x"0c30c3",
   38747 => x"0c30c3",
   38748 => x"0c30c3",
   38749 => x"0c30c3",
   38750 => x"0c30c3",
   38751 => x"0c30c3",
   38752 => x"0c30c3",
   38753 => x"0c30c3",
   38754 => x"0c30c3",
   38755 => x"0c30c3",
   38756 => x"0c30c3",
   38757 => x"0c30c3",
   38758 => x"0c30c3",
   38759 => x"0c30c3",
   38760 => x"0c30c3",
   38761 => x"0c30c3",
   38762 => x"0c30c3",
   38763 => x"0c30c3",
   38764 => x"0c30c3",
   38765 => x"0c30c3",
   38766 => x"0c30c3",
   38767 => x"0c30c3",
   38768 => x"0c30c3",
   38769 => x"0c30c3",
   38770 => x"0c30c3",
   38771 => x"0c30c3",
   38772 => x"0c30c3",
   38773 => x"0c35ff",
   38774 => x"ffffff",
   38775 => x"ffffff",
   38776 => x"ffffff",
   38777 => x"ffffff",
   38778 => x"ffffff",
   38779 => x"ffffff",
   38780 => x"ffffff",
   38781 => x"ffffff",
   38782 => x"ffffff",
   38783 => x"ffffff",
   38784 => x"ffffff",
   38785 => x"ffffff",
   38786 => x"ffffff",
   38787 => x"ffffff",
   38788 => x"ffffff",
   38789 => x"fffa95",
   38790 => x"abffff",
   38791 => x"ffffff",
   38792 => x"ffffff",
   38793 => x"ffffff",
   38794 => x"ffffff",
   38795 => x"ffffff",
   38796 => x"ffffff",
   38797 => x"ffffff",
   38798 => x"ffffff",
   38799 => x"ffffff",
   38800 => x"ffffff",
   38801 => x"fffb8c",
   38802 => x"30c30c",
   38803 => x"30c30c",
   38804 => x"30c30c",
   38805 => x"30c30c",
   38806 => x"30c30c",
   38807 => x"30c30c",
   38808 => x"30c30c",
   38809 => x"30c30c",
   38810 => x"30c30c",
   38811 => x"30c30c",
   38812 => x"30c30c",
   38813 => x"208208",
   38814 => x"208208",
   38815 => x"208208",
   38816 => x"208208",
   38817 => x"208208",
   38818 => x"208208",
   38819 => x"208208",
   38820 => x"208208",
   38821 => x"208208",
   38822 => x"208208",
   38823 => x"208208",
   38824 => x"208208",
   38825 => x"208208",
   38826 => x"208208",
   38827 => x"208208",
   38828 => x"208208",
   38829 => x"208208",
   38830 => x"208208",
   38831 => x"208208",
   38832 => x"208208",
   38833 => x"208208",
   38834 => x"208208",
   38835 => x"208104",
   38836 => x"104104",
   38837 => x"104104",
   38838 => x"104104",
   38839 => x"104104",
   38840 => x"104104",
   38841 => x"104104",
   38842 => x"104104",
   38843 => x"104104",
   38844 => x"104104",
   38845 => x"104104",
   38846 => x"104104",
   38847 => x"104104",
   38848 => x"104104",
   38849 => x"104104",
   38850 => x"104104",
   38851 => x"104104",
   38852 => x"104104",
   38853 => x"104104",
   38854 => x"104104",
   38855 => x"104104",
   38856 => x"104104",
   38857 => x"104104",
   38858 => x"104000",
   38859 => x"000000",
   38860 => x"000000",
   38861 => x"000000",
   38862 => x"000000",
   38863 => x"000000",
   38864 => x"000000",
   38865 => x"000000",
   38866 => x"000000",
   38867 => x"000000",
   38868 => x"000000",
   38869 => x"00057f",
   38870 => x"ffffff",
   38871 => x"ffffff",
   38872 => x"ffffff",
   38873 => x"fff000",
   38874 => x"000abf",
   38875 => x"ffffff",
   38876 => x"ffffff",
   38877 => x"ffffff",
   38878 => x"ffffff",
   38879 => x"ffffff",
   38880 => x"ffffff",
   38881 => x"ffffff",
   38882 => x"ffffff",
   38883 => x"ffffff",
   38884 => x"ffffff",
   38885 => x"ffffff",
   38886 => x"ffffff",
   38887 => x"ffffff",
   38888 => x"ffffff",
   38889 => x"ffffff",
   38890 => x"ffffff",
   38891 => x"ffffff",
   38892 => x"ffffff",
   38893 => x"ffffff",
   38894 => x"ffffff",
   38895 => x"ac30c3",
   38896 => x"0c30c3",
   38897 => x"0c30c3",
   38898 => x"0c30c3",
   38899 => x"0c30c3",
   38900 => x"0c30c3",
   38901 => x"0c30c3",
   38902 => x"0c30c3",
   38903 => x"0c30c3",
   38904 => x"0c30c3",
   38905 => x"0c30c3",
   38906 => x"0c30c3",
   38907 => x"0c30c3",
   38908 => x"0c30c3",
   38909 => x"0c30c3",
   38910 => x"0c30c3",
   38911 => x"0c30c3",
   38912 => x"0c30c3",
   38913 => x"0c30c3",
   38914 => x"0c30c3",
   38915 => x"0c30c3",
   38916 => x"0c30c3",
   38917 => x"0c30c3",
   38918 => x"0c30c3",
   38919 => x"0c30c3",
   38920 => x"0c30c3",
   38921 => x"0c30c3",
   38922 => x"0c30c3",
   38923 => x"0c30c3",
   38924 => x"0c30c3",
   38925 => x"0c30c3",
   38926 => x"0c30c3",
   38927 => x"0c30c3",
   38928 => x"0c30c3",
   38929 => x"0c30c3",
   38930 => x"0c30c3",
   38931 => x"0c30c3",
   38932 => x"0c30c3",
   38933 => x"0d7fff",
   38934 => x"ffffff",
   38935 => x"ffffff",
   38936 => x"ffffff",
   38937 => x"ffffff",
   38938 => x"ffffff",
   38939 => x"ffffff",
   38940 => x"ffffff",
   38941 => x"ffffff",
   38942 => x"ffffff",
   38943 => x"ffffff",
   38944 => x"ffffff",
   38945 => x"ffffff",
   38946 => x"ffffff",
   38947 => x"ffffff",
   38948 => x"ffffff",
   38949 => x"fffa95",
   38950 => x"abffff",
   38951 => x"ffffff",
   38952 => x"ffffff",
   38953 => x"ffffff",
   38954 => x"ffffff",
   38955 => x"ffffff",
   38956 => x"ffffff",
   38957 => x"ffffff",
   38958 => x"ffffff",
   38959 => x"ffffff",
   38960 => x"ffffff",
   38961 => x"fffb8c",
   38962 => x"30c30c",
   38963 => x"30c30c",
   38964 => x"30c30c",
   38965 => x"30c30c",
   38966 => x"30c30c",
   38967 => x"30c30c",
   38968 => x"30c30c",
   38969 => x"30c30c",
   38970 => x"30c30c",
   38971 => x"30c30c",
   38972 => x"30c30c",
   38973 => x"208208",
   38974 => x"208208",
   38975 => x"208208",
   38976 => x"208208",
   38977 => x"208208",
   38978 => x"208208",
   38979 => x"208208",
   38980 => x"208208",
   38981 => x"208208",
   38982 => x"208208",
   38983 => x"208208",
   38984 => x"208208",
   38985 => x"208208",
   38986 => x"208208",
   38987 => x"208208",
   38988 => x"208208",
   38989 => x"208208",
   38990 => x"208208",
   38991 => x"208208",
   38992 => x"208208",
   38993 => x"208208",
   38994 => x"208208",
   38995 => x"208104",
   38996 => x"104104",
   38997 => x"104104",
   38998 => x"104104",
   38999 => x"104104",
   39000 => x"104104",
   39001 => x"104104",
   39002 => x"104104",
   39003 => x"104104",
   39004 => x"104104",
   39005 => x"104104",
   39006 => x"104104",
   39007 => x"104104",
   39008 => x"104104",
   39009 => x"104104",
   39010 => x"104104",
   39011 => x"104104",
   39012 => x"104104",
   39013 => x"104104",
   39014 => x"104104",
   39015 => x"104104",
   39016 => x"104104",
   39017 => x"104104",
   39018 => x"104000",
   39019 => x"000000",
   39020 => x"000000",
   39021 => x"000000",
   39022 => x"000000",
   39023 => x"000000",
   39024 => x"000000",
   39025 => x"000000",
   39026 => x"000000",
   39027 => x"000000",
   39028 => x"000000",
   39029 => x"00057f",
   39030 => x"ffffff",
   39031 => x"ffffff",
   39032 => x"ffffff",
   39033 => x"fea000",
   39034 => x"000abf",
   39035 => x"ffffff",
   39036 => x"ffffff",
   39037 => x"ffffff",
   39038 => x"ffffff",
   39039 => x"ffffff",
   39040 => x"ffffff",
   39041 => x"ffffff",
   39042 => x"ffffff",
   39043 => x"ffffff",
   39044 => x"ffffff",
   39045 => x"ffffff",
   39046 => x"ffffff",
   39047 => x"ffffff",
   39048 => x"ffffff",
   39049 => x"ffffff",
   39050 => x"ffffff",
   39051 => x"ffffff",
   39052 => x"ffffff",
   39053 => x"ffffff",
   39054 => x"ffffff",
   39055 => x"fd70c3",
   39056 => x"0c30c3",
   39057 => x"0c30c3",
   39058 => x"0c30c3",
   39059 => x"0c30c3",
   39060 => x"0c30c3",
   39061 => x"0c30c3",
   39062 => x"0c30c3",
   39063 => x"0c30c3",
   39064 => x"0c30c3",
   39065 => x"0c30c3",
   39066 => x"0c30c3",
   39067 => x"0c30c3",
   39068 => x"0c30c3",
   39069 => x"0c30c3",
   39070 => x"0c30c3",
   39071 => x"0c30c3",
   39072 => x"0c30c3",
   39073 => x"0c30c3",
   39074 => x"0c30c3",
   39075 => x"0c30c3",
   39076 => x"0c30c3",
   39077 => x"0c30c3",
   39078 => x"0c30c3",
   39079 => x"0c30c3",
   39080 => x"0c30c3",
   39081 => x"0c30c3",
   39082 => x"0c30c3",
   39083 => x"0c30c3",
   39084 => x"0c30c3",
   39085 => x"0c30c3",
   39086 => x"0c30c3",
   39087 => x"0c30c3",
   39088 => x"0c30c3",
   39089 => x"0c30c3",
   39090 => x"0c30c3",
   39091 => x"0c30c3",
   39092 => x"0c30c3",
   39093 => x"0ebfff",
   39094 => x"ffffff",
   39095 => x"ffffff",
   39096 => x"ffffff",
   39097 => x"ffffff",
   39098 => x"ffffff",
   39099 => x"ffffff",
   39100 => x"ffffff",
   39101 => x"ffffff",
   39102 => x"ffffff",
   39103 => x"ffffff",
   39104 => x"ffffff",
   39105 => x"ffffff",
   39106 => x"ffffff",
   39107 => x"ffffff",
   39108 => x"ffffff",
   39109 => x"fffa95",
   39110 => x"abffff",
   39111 => x"ffffff",
   39112 => x"ffffff",
   39113 => x"ffffff",
   39114 => x"ffffff",
   39115 => x"ffffff",
   39116 => x"ffffff",
   39117 => x"ffffff",
   39118 => x"ffffff",
   39119 => x"ffffff",
   39120 => x"ffffff",
   39121 => x"fffb8c",
   39122 => x"30c30c",
   39123 => x"30c30c",
   39124 => x"30c30c",
   39125 => x"30c30c",
   39126 => x"30c30c",
   39127 => x"30c30c",
   39128 => x"30c30c",
   39129 => x"30c30c",
   39130 => x"30c30c",
   39131 => x"30c30c",
   39132 => x"30c30c",
   39133 => x"208208",
   39134 => x"208208",
   39135 => x"208208",
   39136 => x"208208",
   39137 => x"208208",
   39138 => x"208208",
   39139 => x"208208",
   39140 => x"208208",
   39141 => x"208208",
   39142 => x"208208",
   39143 => x"208208",
   39144 => x"208208",
   39145 => x"208208",
   39146 => x"208208",
   39147 => x"208208",
   39148 => x"208208",
   39149 => x"208208",
   39150 => x"208208",
   39151 => x"208208",
   39152 => x"208208",
   39153 => x"208208",
   39154 => x"208208",
   39155 => x"208104",
   39156 => x"104104",
   39157 => x"104104",
   39158 => x"104104",
   39159 => x"104104",
   39160 => x"104104",
   39161 => x"104104",
   39162 => x"104104",
   39163 => x"104104",
   39164 => x"104104",
   39165 => x"104104",
   39166 => x"104104",
   39167 => x"104104",
   39168 => x"104104",
   39169 => x"104104",
   39170 => x"104104",
   39171 => x"104104",
   39172 => x"104104",
   39173 => x"104104",
   39174 => x"104104",
   39175 => x"104104",
   39176 => x"104104",
   39177 => x"104104",
   39178 => x"104000",
   39179 => x"000000",
   39180 => x"000000",
   39181 => x"000000",
   39182 => x"000000",
   39183 => x"000000",
   39184 => x"000000",
   39185 => x"000000",
   39186 => x"000000",
   39187 => x"000000",
   39188 => x"000000",
   39189 => x"00057f",
   39190 => x"ffffff",
   39191 => x"ffffff",
   39192 => x"ffffff",
   39193 => x"fea000",
   39194 => x"015fff",
   39195 => x"ffffff",
   39196 => x"ffffff",
   39197 => x"ffffff",
   39198 => x"ffffff",
   39199 => x"ffffff",
   39200 => x"ffffff",
   39201 => x"ffffff",
   39202 => x"ffffff",
   39203 => x"ffffff",
   39204 => x"ffffff",
   39205 => x"ffffff",
   39206 => x"ffffff",
   39207 => x"ffffff",
   39208 => x"ffffff",
   39209 => x"ffffff",
   39210 => x"ffffff",
   39211 => x"ffffff",
   39212 => x"ffffff",
   39213 => x"ffffff",
   39214 => x"ffffff",
   39215 => x"feb5c3",
   39216 => x"0c30c3",
   39217 => x"0c30c3",
   39218 => x"0c30c3",
   39219 => x"0c30c3",
   39220 => x"0c30c3",
   39221 => x"0c30c3",
   39222 => x"0c30c3",
   39223 => x"0c30c3",
   39224 => x"0c30c3",
   39225 => x"0c30c3",
   39226 => x"0c30c3",
   39227 => x"0c30c3",
   39228 => x"0c30c3",
   39229 => x"0c30c3",
   39230 => x"0c30c3",
   39231 => x"0c30c3",
   39232 => x"0c30c3",
   39233 => x"0c30c3",
   39234 => x"0c30c3",
   39235 => x"0c30c3",
   39236 => x"0c30c3",
   39237 => x"0c30c3",
   39238 => x"0c30c3",
   39239 => x"0c30c3",
   39240 => x"0c30c3",
   39241 => x"0c30c3",
   39242 => x"0c30c3",
   39243 => x"0c30c3",
   39244 => x"0c30c3",
   39245 => x"0c30c3",
   39246 => x"0c30c3",
   39247 => x"0c30c3",
   39248 => x"0c30c3",
   39249 => x"0c30c3",
   39250 => x"0c30c3",
   39251 => x"0c30c3",
   39252 => x"0c30c3",
   39253 => x"afffff",
   39254 => x"ffffff",
   39255 => x"ffffff",
   39256 => x"ffffff",
   39257 => x"ffffff",
   39258 => x"ffffff",
   39259 => x"ffffff",
   39260 => x"ffffff",
   39261 => x"ffffff",
   39262 => x"ffffff",
   39263 => x"ffffff",
   39264 => x"ffffff",
   39265 => x"ffffff",
   39266 => x"ffffff",
   39267 => x"ffffff",
   39268 => x"ffffff",
   39269 => x"fffa95",
   39270 => x"abffff",
   39271 => x"ffffff",
   39272 => x"ffffff",
   39273 => x"ffffff",
   39274 => x"ffffff",
   39275 => x"ffffff",
   39276 => x"ffffff",
   39277 => x"ffffff",
   39278 => x"ffffff",
   39279 => x"ffffff",
   39280 => x"ffffff",
   39281 => x"fffb8c",
   39282 => x"30c30c",
   39283 => x"30c30c",
   39284 => x"30c30c",
   39285 => x"30c30c",
   39286 => x"30c30c",
   39287 => x"30c30c",
   39288 => x"30c30c",
   39289 => x"30c30c",
   39290 => x"30c30c",
   39291 => x"30c30c",
   39292 => x"30c30c",
   39293 => x"208208",
   39294 => x"208208",
   39295 => x"208208",
   39296 => x"208208",
   39297 => x"208208",
   39298 => x"208208",
   39299 => x"208208",
   39300 => x"208208",
   39301 => x"208208",
   39302 => x"208208",
   39303 => x"208208",
   39304 => x"208208",
   39305 => x"208208",
   39306 => x"208208",
   39307 => x"208208",
   39308 => x"208208",
   39309 => x"208208",
   39310 => x"208208",
   39311 => x"208208",
   39312 => x"208208",
   39313 => x"208208",
   39314 => x"208208",
   39315 => x"208104",
   39316 => x"104104",
   39317 => x"104104",
   39318 => x"104104",
   39319 => x"104104",
   39320 => x"104104",
   39321 => x"104104",
   39322 => x"104104",
   39323 => x"104104",
   39324 => x"104104",
   39325 => x"104104",
   39326 => x"104104",
   39327 => x"104104",
   39328 => x"104104",
   39329 => x"104104",
   39330 => x"104104",
   39331 => x"104104",
   39332 => x"104104",
   39333 => x"104104",
   39334 => x"104104",
   39335 => x"104104",
   39336 => x"104104",
   39337 => x"104104",
   39338 => x"104000",
   39339 => x"000000",
   39340 => x"000000",
   39341 => x"000000",
   39342 => x"000000",
   39343 => x"000000",
   39344 => x"000000",
   39345 => x"000000",
   39346 => x"000000",
   39347 => x"000000",
   39348 => x"000000",
   39349 => x"00057f",
   39350 => x"ffffff",
   39351 => x"ffffff",
   39352 => x"ffffff",
   39353 => x"fea000",
   39354 => x"015fff",
   39355 => x"ffffff",
   39356 => x"ffffff",
   39357 => x"feaaaa",
   39358 => x"aaaaaa",
   39359 => x"aaaaaa",
   39360 => x"ffffff",
   39361 => x"ffffff",
   39362 => x"ffffff",
   39363 => x"ffffff",
   39364 => x"ffffff",
   39365 => x"ffffff",
   39366 => x"ffffff",
   39367 => x"ffffff",
   39368 => x"ffffff",
   39369 => x"ffffff",
   39370 => x"ffffff",
   39371 => x"ffffff",
   39372 => x"ffffff",
   39373 => x"ffffff",
   39374 => x"ffffff",
   39375 => x"fffad7",
   39376 => x"0c30c3",
   39377 => x"0c30c3",
   39378 => x"0c30c3",
   39379 => x"0c30c3",
   39380 => x"0c30c3",
   39381 => x"0c30c3",
   39382 => x"0c30c3",
   39383 => x"0c30c3",
   39384 => x"0c30c3",
   39385 => x"0c30c3",
   39386 => x"0c30c3",
   39387 => x"0c30c3",
   39388 => x"0c30c3",
   39389 => x"0c30c3",
   39390 => x"0c30c3",
   39391 => x"0c30c3",
   39392 => x"0c30c3",
   39393 => x"0c30c3",
   39394 => x"0c30c3",
   39395 => x"0c30c3",
   39396 => x"0c30c3",
   39397 => x"0c30c3",
   39398 => x"0c30c3",
   39399 => x"0c30c3",
   39400 => x"0c30c3",
   39401 => x"0c30c3",
   39402 => x"0c30c3",
   39403 => x"0c30c3",
   39404 => x"0c30c3",
   39405 => x"0c30c3",
   39406 => x"0c30c3",
   39407 => x"0c30c3",
   39408 => x"0c30c3",
   39409 => x"0c30c3",
   39410 => x"0c30c3",
   39411 => x"0c30c3",
   39412 => x"0c30d7",
   39413 => x"ffffff",
   39414 => x"ffffff",
   39415 => x"ffffff",
   39416 => x"ffffff",
   39417 => x"ffffff",
   39418 => x"ffffff",
   39419 => x"ffffff",
   39420 => x"ffffff",
   39421 => x"ffffff",
   39422 => x"ffffff",
   39423 => x"ffffff",
   39424 => x"ffffff",
   39425 => x"ffffff",
   39426 => x"ffffff",
   39427 => x"ffffff",
   39428 => x"ffffff",
   39429 => x"fffa95",
   39430 => x"abffff",
   39431 => x"ffffff",
   39432 => x"ffffff",
   39433 => x"ffffff",
   39434 => x"ffffff",
   39435 => x"ffffff",
   39436 => x"ffffff",
   39437 => x"ffffff",
   39438 => x"ffffff",
   39439 => x"ffffff",
   39440 => x"ffffff",
   39441 => x"fffb8c",
   39442 => x"30c30c",
   39443 => x"30c30c",
   39444 => x"30c30c",
   39445 => x"30c30c",
   39446 => x"30c30c",
   39447 => x"30c30c",
   39448 => x"30c30c",
   39449 => x"30c30c",
   39450 => x"30c30c",
   39451 => x"30c30c",
   39452 => x"30c30c",
   39453 => x"208208",
   39454 => x"208208",
   39455 => x"208208",
   39456 => x"208208",
   39457 => x"208208",
   39458 => x"208208",
   39459 => x"208208",
   39460 => x"208208",
   39461 => x"208208",
   39462 => x"208208",
   39463 => x"208208",
   39464 => x"208208",
   39465 => x"208208",
   39466 => x"208208",
   39467 => x"208208",
   39468 => x"208208",
   39469 => x"208208",
   39470 => x"208208",
   39471 => x"208208",
   39472 => x"208208",
   39473 => x"208208",
   39474 => x"208208",
   39475 => x"208104",
   39476 => x"104104",
   39477 => x"104104",
   39478 => x"104104",
   39479 => x"104104",
   39480 => x"104104",
   39481 => x"104104",
   39482 => x"104104",
   39483 => x"104104",
   39484 => x"104104",
   39485 => x"104104",
   39486 => x"104104",
   39487 => x"104104",
   39488 => x"104104",
   39489 => x"104104",
   39490 => x"104104",
   39491 => x"104104",
   39492 => x"104104",
   39493 => x"104104",
   39494 => x"104104",
   39495 => x"104104",
   39496 => x"104104",
   39497 => x"104104",
   39498 => x"104000",
   39499 => x"000000",
   39500 => x"000000",
   39501 => x"000000",
   39502 => x"000000",
   39503 => x"000000",
   39504 => x"000000",
   39505 => x"000000",
   39506 => x"000000",
   39507 => x"000000",
   39508 => x"000000",
   39509 => x"00057f",
   39510 => x"ffffff",
   39511 => x"ffffff",
   39512 => x"ffffff",
   39513 => x"fea000",
   39514 => x"015fff",
   39515 => x"ffffff",
   39516 => x"ffffff",
   39517 => x"fd5015",
   39518 => x"555555",
   39519 => x"555555",
   39520 => x"ffffff",
   39521 => x"ffffff",
   39522 => x"ffffff",
   39523 => x"ffffff",
   39524 => x"ffffff",
   39525 => x"ffffff",
   39526 => x"ffffff",
   39527 => x"ffffff",
   39528 => x"ffffff",
   39529 => x"ffffff",
   39530 => x"ffffff",
   39531 => x"ffffff",
   39532 => x"ffffff",
   39533 => x"ffffff",
   39534 => x"ffffff",
   39535 => x"ffffeb",
   39536 => x"0c30c3",
   39537 => x"0c30c3",
   39538 => x"0c30c3",
   39539 => x"0c30c3",
   39540 => x"0c30c3",
   39541 => x"0c30c3",
   39542 => x"0c30c3",
   39543 => x"0c30c3",
   39544 => x"0c30c3",
   39545 => x"0c30c3",
   39546 => x"0c30c3",
   39547 => x"0c30c3",
   39548 => x"0c30c3",
   39549 => x"0c30c3",
   39550 => x"0c30c3",
   39551 => x"0c30c3",
   39552 => x"0c30c3",
   39553 => x"0c30c3",
   39554 => x"0c30c3",
   39555 => x"0c30c3",
   39556 => x"0c30c3",
   39557 => x"0c30c3",
   39558 => x"0c30c3",
   39559 => x"0c30c3",
   39560 => x"0c30c3",
   39561 => x"0c30c3",
   39562 => x"0c30c3",
   39563 => x"0c30c3",
   39564 => x"0c30c3",
   39565 => x"0c30c3",
   39566 => x"0c30c3",
   39567 => x"0c30c3",
   39568 => x"0c30c3",
   39569 => x"0c30c3",
   39570 => x"0c30c3",
   39571 => x"0c30c3",
   39572 => x"0c35eb",
   39573 => x"ffffff",
   39574 => x"ffffff",
   39575 => x"ffffff",
   39576 => x"ffffff",
   39577 => x"ffffff",
   39578 => x"ffffff",
   39579 => x"ffffff",
   39580 => x"ffffff",
   39581 => x"ffffff",
   39582 => x"ffffff",
   39583 => x"ffffff",
   39584 => x"ffffff",
   39585 => x"ffffff",
   39586 => x"ffffff",
   39587 => x"ffffff",
   39588 => x"ffffff",
   39589 => x"fffa95",
   39590 => x"abffff",
   39591 => x"ffffff",
   39592 => x"ffffff",
   39593 => x"ffffff",
   39594 => x"ffffff",
   39595 => x"ffffff",
   39596 => x"ffffff",
   39597 => x"ffffff",
   39598 => x"ffffff",
   39599 => x"ffffff",
   39600 => x"ffffff",
   39601 => x"fffb8c",
   39602 => x"30c30c",
   39603 => x"30c30c",
   39604 => x"30c30c",
   39605 => x"30c30c",
   39606 => x"30c30c",
   39607 => x"30c30c",
   39608 => x"30c30c",
   39609 => x"30c30c",
   39610 => x"30c30c",
   39611 => x"30c30c",
   39612 => x"30c30c",
   39613 => x"208208",
   39614 => x"208208",
   39615 => x"208208",
   39616 => x"208208",
   39617 => x"208208",
   39618 => x"208208",
   39619 => x"208208",
   39620 => x"208208",
   39621 => x"208208",
   39622 => x"208208",
   39623 => x"208208",
   39624 => x"208208",
   39625 => x"208208",
   39626 => x"208208",
   39627 => x"208208",
   39628 => x"208208",
   39629 => x"208208",
   39630 => x"208208",
   39631 => x"208208",
   39632 => x"208208",
   39633 => x"208208",
   39634 => x"208208",
   39635 => x"208104",
   39636 => x"104104",
   39637 => x"104104",
   39638 => x"104104",
   39639 => x"104104",
   39640 => x"104104",
   39641 => x"104104",
   39642 => x"104104",
   39643 => x"104104",
   39644 => x"104104",
   39645 => x"104104",
   39646 => x"104104",
   39647 => x"104104",
   39648 => x"104104",
   39649 => x"104104",
   39650 => x"104104",
   39651 => x"104104",
   39652 => x"104104",
   39653 => x"104104",
   39654 => x"104104",
   39655 => x"104104",
   39656 => x"104104",
   39657 => x"104104",
   39658 => x"104000",
   39659 => x"000000",
   39660 => x"000000",
   39661 => x"000000",
   39662 => x"000000",
   39663 => x"000000",
   39664 => x"000000",
   39665 => x"000000",
   39666 => x"000000",
   39667 => x"000000",
   39668 => x"000000",
   39669 => x"00057f",
   39670 => x"ffffff",
   39671 => x"ffffff",
   39672 => x"ffffff",
   39673 => x"fea000",
   39674 => x"015fff",
   39675 => x"ffffff",
   39676 => x"ffffff",
   39677 => x"fd5000",
   39678 => x"000000",
   39679 => x"000000",
   39680 => x"ffffff",
   39681 => x"ffffff",
   39682 => x"ffffff",
   39683 => x"ffffff",
   39684 => x"ffffff",
   39685 => x"ffffff",
   39686 => x"ffffff",
   39687 => x"ffffff",
   39688 => x"ffffff",
   39689 => x"ffffff",
   39690 => x"ffffff",
   39691 => x"ffffff",
   39692 => x"ffffff",
   39693 => x"ffffff",
   39694 => x"ffffff",
   39695 => x"ffffff",
   39696 => x"5c30c3",
   39697 => x"0c30c3",
   39698 => x"0c30c3",
   39699 => x"0c30c3",
   39700 => x"0c30c3",
   39701 => x"0c30c3",
   39702 => x"0c30c3",
   39703 => x"0c30c3",
   39704 => x"0c30c3",
   39705 => x"0c30c3",
   39706 => x"0c30c3",
   39707 => x"0c30c3",
   39708 => x"0c30c3",
   39709 => x"0c30c3",
   39710 => x"0c30c3",
   39711 => x"0c30c3",
   39712 => x"0c30c3",
   39713 => x"0c30c3",
   39714 => x"0c30c3",
   39715 => x"0c30c3",
   39716 => x"0c30c3",
   39717 => x"0c30c3",
   39718 => x"0c30c3",
   39719 => x"0c30c3",
   39720 => x"0c30c3",
   39721 => x"0c30c3",
   39722 => x"0c30c3",
   39723 => x"0c30c3",
   39724 => x"0c30c3",
   39725 => x"0c30c3",
   39726 => x"0c30c3",
   39727 => x"0c30c3",
   39728 => x"0c30c3",
   39729 => x"0c30c3",
   39730 => x"0c30c3",
   39731 => x"0c30c3",
   39732 => x"0c3aff",
   39733 => x"ffffff",
   39734 => x"ffffff",
   39735 => x"ffffff",
   39736 => x"ffffff",
   39737 => x"ffffff",
   39738 => x"ffffff",
   39739 => x"ffffff",
   39740 => x"ffffff",
   39741 => x"ffffff",
   39742 => x"ffffff",
   39743 => x"ffffff",
   39744 => x"ffffff",
   39745 => x"ffffff",
   39746 => x"ffffff",
   39747 => x"ffffff",
   39748 => x"ffffff",
   39749 => x"fffa95",
   39750 => x"abffff",
   39751 => x"ffffff",
   39752 => x"ffffff",
   39753 => x"ffffff",
   39754 => x"ffffff",
   39755 => x"ffffff",
   39756 => x"ffffff",
   39757 => x"ffffff",
   39758 => x"ffffff",
   39759 => x"ffffff",
   39760 => x"ffffff",
   39761 => x"fffb8c",
   39762 => x"30c30c",
   39763 => x"30c30c",
   39764 => x"30c30c",
   39765 => x"30c30c",
   39766 => x"30c30c",
   39767 => x"30c30c",
   39768 => x"30c30c",
   39769 => x"30c30c",
   39770 => x"30c30c",
   39771 => x"30c30c",
   39772 => x"30c30c",
   39773 => x"208208",
   39774 => x"208208",
   39775 => x"208208",
   39776 => x"208208",
   39777 => x"208208",
   39778 => x"208208",
   39779 => x"208208",
   39780 => x"208208",
   39781 => x"208208",
   39782 => x"208208",
   39783 => x"208208",
   39784 => x"208208",
   39785 => x"208208",
   39786 => x"208208",
   39787 => x"208208",
   39788 => x"208208",
   39789 => x"208208",
   39790 => x"208208",
   39791 => x"208208",
   39792 => x"208208",
   39793 => x"208208",
   39794 => x"208208",
   39795 => x"208104",
   39796 => x"104104",
   39797 => x"104104",
   39798 => x"104104",
   39799 => x"104104",
   39800 => x"104104",
   39801 => x"104104",
   39802 => x"104104",
   39803 => x"104104",
   39804 => x"104104",
   39805 => x"104104",
   39806 => x"104104",
   39807 => x"104104",
   39808 => x"104104",
   39809 => x"104104",
   39810 => x"104104",
   39811 => x"104104",
   39812 => x"104104",
   39813 => x"104104",
   39814 => x"104104",
   39815 => x"104104",
   39816 => x"104104",
   39817 => x"104104",
   39818 => x"104000",
   39819 => x"000000",
   39820 => x"000000",
   39821 => x"000000",
   39822 => x"000000",
   39823 => x"000000",
   39824 => x"000000",
   39825 => x"000000",
   39826 => x"000000",
   39827 => x"000000",
   39828 => x"000000",
   39829 => x"00057f",
   39830 => x"ffffff",
   39831 => x"ffffff",
   39832 => x"ffffff",
   39833 => x"fea000",
   39834 => x"015fff",
   39835 => x"ffffff",
   39836 => x"ffffff",
   39837 => x"fd5000",
   39838 => x"000000",
   39839 => x"000000",
   39840 => x"ffffff",
   39841 => x"ffffff",
   39842 => x"ffffff",
   39843 => x"ffffff",
   39844 => x"ffffff",
   39845 => x"ffffff",
   39846 => x"ffffff",
   39847 => x"ffffff",
   39848 => x"ffffff",
   39849 => x"ffffff",
   39850 => x"ffffff",
   39851 => x"ffffff",
   39852 => x"ffffff",
   39853 => x"ffffff",
   39854 => x"ffffff",
   39855 => x"ffffff",
   39856 => x"ad70c3",
   39857 => x"0c30c3",
   39858 => x"0c30c3",
   39859 => x"0c30c3",
   39860 => x"0c30c3",
   39861 => x"0c30c3",
   39862 => x"0c30c3",
   39863 => x"0c30c3",
   39864 => x"0c30c3",
   39865 => x"0c30c3",
   39866 => x"0c30c3",
   39867 => x"0c30c3",
   39868 => x"0c30c3",
   39869 => x"0c30c3",
   39870 => x"0c30c3",
   39871 => x"0c30c3",
   39872 => x"0c30c3",
   39873 => x"0c30c3",
   39874 => x"0c30c3",
   39875 => x"0c30c3",
   39876 => x"0c30c3",
   39877 => x"0c30c3",
   39878 => x"0c30c3",
   39879 => x"0c30c3",
   39880 => x"0c30c3",
   39881 => x"0c30c3",
   39882 => x"0c30c3",
   39883 => x"0c30c3",
   39884 => x"0c30c3",
   39885 => x"0c30c3",
   39886 => x"0c30c3",
   39887 => x"0c30c3",
   39888 => x"0c30c3",
   39889 => x"0c30c3",
   39890 => x"0c30c3",
   39891 => x"0c30c3",
   39892 => x"0d7fff",
   39893 => x"ffffff",
   39894 => x"ffffff",
   39895 => x"ffffff",
   39896 => x"ffffff",
   39897 => x"ffffff",
   39898 => x"ffffff",
   39899 => x"ffffff",
   39900 => x"ffffff",
   39901 => x"ffffff",
   39902 => x"ffffff",
   39903 => x"ffffff",
   39904 => x"ffffff",
   39905 => x"ffffff",
   39906 => x"ffffff",
   39907 => x"ffffff",
   39908 => x"ffffff",
   39909 => x"fffa95",
   39910 => x"abffff",
   39911 => x"ffffff",
   39912 => x"ffffff",
   39913 => x"ffffff",
   39914 => x"ffffff",
   39915 => x"ffffff",
   39916 => x"ffffff",
   39917 => x"ffffff",
   39918 => x"ffffff",
   39919 => x"ffffff",
   39920 => x"ffffff",
   39921 => x"fffb8c",
   39922 => x"30c30c",
   39923 => x"30c30c",
   39924 => x"30c30c",
   39925 => x"30c30c",
   39926 => x"30c30c",
   39927 => x"30c30c",
   39928 => x"30c30c",
   39929 => x"30c30c",
   39930 => x"30c30c",
   39931 => x"30c30c",
   39932 => x"30c30c",
   39933 => x"208208",
   39934 => x"208208",
   39935 => x"208208",
   39936 => x"208208",
   39937 => x"208208",
   39938 => x"208208",
   39939 => x"208208",
   39940 => x"208208",
   39941 => x"208208",
   39942 => x"208208",
   39943 => x"208208",
   39944 => x"208208",
   39945 => x"208208",
   39946 => x"208208",
   39947 => x"208208",
   39948 => x"208208",
   39949 => x"208208",
   39950 => x"208208",
   39951 => x"208208",
   39952 => x"208208",
   39953 => x"208208",
   39954 => x"208208",
   39955 => x"208104",
   39956 => x"104104",
   39957 => x"104104",
   39958 => x"104104",
   39959 => x"104104",
   39960 => x"104104",
   39961 => x"104104",
   39962 => x"104104",
   39963 => x"104104",
   39964 => x"104104",
   39965 => x"104104",
   39966 => x"104104",
   39967 => x"104104",
   39968 => x"104104",
   39969 => x"104104",
   39970 => x"104104",
   39971 => x"104104",
   39972 => x"104104",
   39973 => x"104104",
   39974 => x"104104",
   39975 => x"104104",
   39976 => x"104104",
   39977 => x"104104",
   39978 => x"104000",
   39979 => x"000000",
   39980 => x"000000",
   39981 => x"000000",
   39982 => x"000000",
   39983 => x"000000",
   39984 => x"000000",
   39985 => x"000000",
   39986 => x"000000",
   39987 => x"000000",
   39988 => x"000000",
   39989 => x"00057f",
   39990 => x"ffffff",
   39991 => x"ffffff",
   39992 => x"ffffff",
   39993 => x"fea000",
   39994 => x"000fff",
   39995 => x"ffffff",
   39996 => x"ffffff",
   39997 => x"feaaaa",
   39998 => x"aaaaaa",
   39999 => x"000000",
   40000 => x"ffffff",
   40001 => x"ffffff",
   40002 => x"ffffff",
   40003 => x"ffffff",
   40004 => x"ffffff",
   40005 => x"ffffff",
   40006 => x"ffffff",
   40007 => x"ffffff",
   40008 => x"ffffff",
   40009 => x"ffffff",
   40010 => x"ffffff",
   40011 => x"ffffff",
   40012 => x"ffffff",
   40013 => x"ffffff",
   40014 => x"ffffff",
   40015 => x"ffffff",
   40016 => x"feb5c3",
   40017 => x"0c30c3",
   40018 => x"0c30c3",
   40019 => x"0c30c3",
   40020 => x"0c30c3",
   40021 => x"0c30c3",
   40022 => x"0c30c3",
   40023 => x"0c30c3",
   40024 => x"0c30c3",
   40025 => x"0c30c3",
   40026 => x"0c30c3",
   40027 => x"0c30c3",
   40028 => x"0c30c3",
   40029 => x"0c30c3",
   40030 => x"0c30c3",
   40031 => x"0c30c3",
   40032 => x"0c30c3",
   40033 => x"0c30c3",
   40034 => x"0c30c3",
   40035 => x"0c30c3",
   40036 => x"0c30c3",
   40037 => x"0c30c3",
   40038 => x"0c30c3",
   40039 => x"0c30c3",
   40040 => x"0c30c3",
   40041 => x"0c30c3",
   40042 => x"0c30c3",
   40043 => x"0c30c3",
   40044 => x"0c30c3",
   40045 => x"0c30c3",
   40046 => x"0c30c3",
   40047 => x"0c30c3",
   40048 => x"0c30c3",
   40049 => x"0c30c3",
   40050 => x"0c30c3",
   40051 => x"0c30c3",
   40052 => x"5fffff",
   40053 => x"ffffff",
   40054 => x"ffffff",
   40055 => x"ffffff",
   40056 => x"ffffff",
   40057 => x"ffffff",
   40058 => x"ffffff",
   40059 => x"ffffff",
   40060 => x"ffffff",
   40061 => x"ffffff",
   40062 => x"ffffff",
   40063 => x"ffffff",
   40064 => x"ffffff",
   40065 => x"ffffff",
   40066 => x"ffffff",
   40067 => x"ffffff",
   40068 => x"ffffff",
   40069 => x"fffa95",
   40070 => x"abffff",
   40071 => x"ffffff",
   40072 => x"ffffff",
   40073 => x"ffffff",
   40074 => x"ffffff",
   40075 => x"ffffff",
   40076 => x"ffffff",
   40077 => x"ffffff",
   40078 => x"ffffff",
   40079 => x"ffffff",
   40080 => x"ffffff",
   40081 => x"fffb8c",
   40082 => x"30c30c",
   40083 => x"30c30c",
   40084 => x"30c30c",
   40085 => x"30c30c",
   40086 => x"30c30c",
   40087 => x"30c30c",
   40088 => x"30c30c",
   40089 => x"30c30c",
   40090 => x"30c30c",
   40091 => x"30c30c",
   40092 => x"30c30c",
   40093 => x"208208",
   40094 => x"208208",
   40095 => x"208208",
   40096 => x"208208",
   40097 => x"208208",
   40098 => x"208208",
   40099 => x"208208",
   40100 => x"208208",
   40101 => x"208208",
   40102 => x"208208",
   40103 => x"208208",
   40104 => x"208208",
   40105 => x"208208",
   40106 => x"208208",
   40107 => x"208208",
   40108 => x"208208",
   40109 => x"208208",
   40110 => x"208208",
   40111 => x"208208",
   40112 => x"208208",
   40113 => x"208208",
   40114 => x"208208",
   40115 => x"208104",
   40116 => x"104104",
   40117 => x"104104",
   40118 => x"104104",
   40119 => x"104104",
   40120 => x"104104",
   40121 => x"104104",
   40122 => x"104104",
   40123 => x"104104",
   40124 => x"104104",
   40125 => x"104104",
   40126 => x"104104",
   40127 => x"104104",
   40128 => x"104104",
   40129 => x"104104",
   40130 => x"104104",
   40131 => x"104104",
   40132 => x"104104",
   40133 => x"104104",
   40134 => x"104104",
   40135 => x"104104",
   40136 => x"104104",
   40137 => x"104104",
   40138 => x"104000",
   40139 => x"000000",
   40140 => x"000000",
   40141 => x"000000",
   40142 => x"000000",
   40143 => x"000000",
   40144 => x"000000",
   40145 => x"000000",
   40146 => x"000000",
   40147 => x"000000",
   40148 => x"000000",
   40149 => x"00057f",
   40150 => x"ffffff",
   40151 => x"ffffff",
   40152 => x"ffffff",
   40153 => x"fff000",
   40154 => x"000abf",
   40155 => x"ffffff",
   40156 => x"ffffff",
   40157 => x"ffffff",
   40158 => x"ffffff",
   40159 => x"000000",
   40160 => x"ffffff",
   40161 => x"ffffff",
   40162 => x"ffffff",
   40163 => x"ffffff",
   40164 => x"ffffff",
   40165 => x"ffffff",
   40166 => x"ffffff",
   40167 => x"ffffff",
   40168 => x"ffffff",
   40169 => x"ffffff",
   40170 => x"ffffff",
   40171 => x"ffffff",
   40172 => x"ffffff",
   40173 => x"ffffff",
   40174 => x"ffffff",
   40175 => x"ffffff",
   40176 => x"fffac3",
   40177 => x"0c30c3",
   40178 => x"0c30c3",
   40179 => x"0c30c3",
   40180 => x"0c30c3",
   40181 => x"0c30c3",
   40182 => x"0c30c3",
   40183 => x"0c30c3",
   40184 => x"0c30c3",
   40185 => x"0c30c3",
   40186 => x"0c30c3",
   40187 => x"0c30c3",
   40188 => x"0c30c3",
   40189 => x"0c30c3",
   40190 => x"0c30c3",
   40191 => x"0c30c3",
   40192 => x"0c30c3",
   40193 => x"0c30c3",
   40194 => x"0c30c3",
   40195 => x"0c30c3",
   40196 => x"0c30c3",
   40197 => x"0c30c3",
   40198 => x"0c30c3",
   40199 => x"0c30c3",
   40200 => x"0c30c3",
   40201 => x"0c30c3",
   40202 => x"0c30c3",
   40203 => x"0c30c3",
   40204 => x"0c30c3",
   40205 => x"0c30c3",
   40206 => x"0c30c3",
   40207 => x"0c30c3",
   40208 => x"0c30c3",
   40209 => x"0c30c3",
   40210 => x"0c30c3",
   40211 => x"0c30d7",
   40212 => x"afffff",
   40213 => x"ffffff",
   40214 => x"ffffff",
   40215 => x"ffffff",
   40216 => x"ffffff",
   40217 => x"ffffff",
   40218 => x"ffffff",
   40219 => x"ffffff",
   40220 => x"ffffff",
   40221 => x"ffffff",
   40222 => x"ffffff",
   40223 => x"ffffff",
   40224 => x"ffffff",
   40225 => x"ffffff",
   40226 => x"ffffff",
   40227 => x"ffffff",
   40228 => x"ffffff",
   40229 => x"fffa95",
   40230 => x"abffff",
   40231 => x"ffffff",
   40232 => x"ffffff",
   40233 => x"ffffff",
   40234 => x"ffffff",
   40235 => x"ffffff",
   40236 => x"ffffff",
   40237 => x"ffffff",
   40238 => x"ffffff",
   40239 => x"ffffff",
   40240 => x"ffffff",
   40241 => x"fffb8c",
   40242 => x"30c30c",
   40243 => x"30c30c",
   40244 => x"30c30c",
   40245 => x"30c30c",
   40246 => x"30c30c",
   40247 => x"30c30c",
   40248 => x"30c30c",
   40249 => x"30c30c",
   40250 => x"30c30c",
   40251 => x"30c30c",
   40252 => x"30c30c",
   40253 => x"208208",
   40254 => x"208208",
   40255 => x"208208",
   40256 => x"208208",
   40257 => x"208208",
   40258 => x"208208",
   40259 => x"208208",
   40260 => x"208208",
   40261 => x"208208",
   40262 => x"208208",
   40263 => x"208208",
   40264 => x"208208",
   40265 => x"208208",
   40266 => x"208208",
   40267 => x"208208",
   40268 => x"208208",
   40269 => x"208208",
   40270 => x"208208",
   40271 => x"208208",
   40272 => x"208208",
   40273 => x"208208",
   40274 => x"208208",
   40275 => x"208104",
   40276 => x"104104",
   40277 => x"104104",
   40278 => x"104104",
   40279 => x"104104",
   40280 => x"104104",
   40281 => x"104104",
   40282 => x"104104",
   40283 => x"104104",
   40284 => x"104104",
   40285 => x"104104",
   40286 => x"104104",
   40287 => x"104104",
   40288 => x"104104",
   40289 => x"104104",
   40290 => x"104104",
   40291 => x"104104",
   40292 => x"104104",
   40293 => x"104104",
   40294 => x"104104",
   40295 => x"104104",
   40296 => x"104104",
   40297 => x"104104",
   40298 => x"104000",
   40299 => x"000000",
   40300 => x"000000",
   40301 => x"000000",
   40302 => x"000000",
   40303 => x"000000",
   40304 => x"000000",
   40305 => x"000000",
   40306 => x"000000",
   40307 => x"000000",
   40308 => x"000000",
   40309 => x"00057f",
   40310 => x"ffffff",
   40311 => x"ffffff",
   40312 => x"ffffff",
   40313 => x"fff540",
   40314 => x"000abf",
   40315 => x"ffffff",
   40316 => x"ffffff",
   40317 => x"ffffff",
   40318 => x"ffffff",
   40319 => x"000000",
   40320 => x"ffffff",
   40321 => x"ffffff",
   40322 => x"ffffff",
   40323 => x"ffffff",
   40324 => x"ffffff",
   40325 => x"ffffff",
   40326 => x"ffffff",
   40327 => x"ffffff",
   40328 => x"ffffff",
   40329 => x"ffffff",
   40330 => x"ffffff",
   40331 => x"ffffff",
   40332 => x"ffffff",
   40333 => x"ffffff",
   40334 => x"ffffff",
   40335 => x"ffffff",
   40336 => x"ffffeb",
   40337 => x"0c30c3",
   40338 => x"0c30c3",
   40339 => x"0c30c3",
   40340 => x"0c30c3",
   40341 => x"0c30c3",
   40342 => x"0c30c3",
   40343 => x"0c30c3",
   40344 => x"0c30c3",
   40345 => x"0c30c3",
   40346 => x"0c30c3",
   40347 => x"0c30c3",
   40348 => x"0c30c3",
   40349 => x"0c30c3",
   40350 => x"0c30c3",
   40351 => x"0c30c3",
   40352 => x"0c30c3",
   40353 => x"0c30c3",
   40354 => x"0c30c3",
   40355 => x"0c30c3",
   40356 => x"0c30c3",
   40357 => x"0c30c3",
   40358 => x"0c30c3",
   40359 => x"0c30c3",
   40360 => x"0c30c3",
   40361 => x"0c30c3",
   40362 => x"0c30c3",
   40363 => x"0c30c3",
   40364 => x"0c30c3",
   40365 => x"0c30c3",
   40366 => x"0c30c3",
   40367 => x"0c30c3",
   40368 => x"0c30c3",
   40369 => x"0c30c3",
   40370 => x"0c30c3",
   40371 => x"0c35eb",
   40372 => x"ffffff",
   40373 => x"ffffff",
   40374 => x"ffffff",
   40375 => x"ffffff",
   40376 => x"ffffff",
   40377 => x"ffffff",
   40378 => x"ffffff",
   40379 => x"ffffff",
   40380 => x"ffffff",
   40381 => x"ffffff",
   40382 => x"ffffff",
   40383 => x"ffffff",
   40384 => x"ffffff",
   40385 => x"ffffff",
   40386 => x"ffffff",
   40387 => x"ffffff",
   40388 => x"ffffff",
   40389 => x"fffa95",
   40390 => x"abffff",
   40391 => x"ffffff",
   40392 => x"ffffff",
   40393 => x"ffffff",
   40394 => x"ffffff",
   40395 => x"ffffff",
   40396 => x"ffffff",
   40397 => x"ffffff",
   40398 => x"ffffff",
   40399 => x"ffffff",
   40400 => x"ffffff",
   40401 => x"fffb8c",
   40402 => x"30c30c",
   40403 => x"30c30c",
   40404 => x"30c30c",
   40405 => x"30c30c",
   40406 => x"30c30c",
   40407 => x"30c30c",
   40408 => x"30c30c",
   40409 => x"30c30c",
   40410 => x"30c30c",
   40411 => x"30c30c",
   40412 => x"30c30c",
   40413 => x"208208",
   40414 => x"208208",
   40415 => x"208208",
   40416 => x"208208",
   40417 => x"208208",
   40418 => x"208208",
   40419 => x"208208",
   40420 => x"208208",
   40421 => x"208208",
   40422 => x"208208",
   40423 => x"208208",
   40424 => x"208208",
   40425 => x"208208",
   40426 => x"208208",
   40427 => x"208208",
   40428 => x"208208",
   40429 => x"208208",
   40430 => x"208208",
   40431 => x"208208",
   40432 => x"208208",
   40433 => x"208208",
   40434 => x"208208",
   40435 => x"208104",
   40436 => x"104104",
   40437 => x"104104",
   40438 => x"104104",
   40439 => x"104104",
   40440 => x"104104",
   40441 => x"104104",
   40442 => x"104104",
   40443 => x"104104",
   40444 => x"104104",
   40445 => x"104104",
   40446 => x"104104",
   40447 => x"104104",
   40448 => x"104104",
   40449 => x"104104",
   40450 => x"104104",
   40451 => x"104104",
   40452 => x"104104",
   40453 => x"104104",
   40454 => x"104104",
   40455 => x"104104",
   40456 => x"104104",
   40457 => x"104104",
   40458 => x"104000",
   40459 => x"000000",
   40460 => x"000000",
   40461 => x"000000",
   40462 => x"000000",
   40463 => x"000000",
   40464 => x"000000",
   40465 => x"000000",
   40466 => x"000000",
   40467 => x"000000",
   40468 => x"000000",
   40469 => x"00057f",
   40470 => x"ffffff",
   40471 => x"ffffff",
   40472 => x"ffffff",
   40473 => x"fff540",
   40474 => x"00057f",
   40475 => x"ffffff",
   40476 => x"ffffff",
   40477 => x"ffffff",
   40478 => x"ffffff",
   40479 => x"000000",
   40480 => x"ffffff",
   40481 => x"ffffff",
   40482 => x"ffffff",
   40483 => x"ffffff",
   40484 => x"ffffff",
   40485 => x"ffffff",
   40486 => x"ffffff",
   40487 => x"ffffff",
   40488 => x"ffffff",
   40489 => x"ffffff",
   40490 => x"ffffff",
   40491 => x"ffffff",
   40492 => x"ffffff",
   40493 => x"ffffff",
   40494 => x"ffffff",
   40495 => x"ffffff",
   40496 => x"ffffff",
   40497 => x"ac30c3",
   40498 => x"0c30c3",
   40499 => x"0c30c3",
   40500 => x"0c30c3",
   40501 => x"0c30c3",
   40502 => x"0c30c3",
   40503 => x"0c30c3",
   40504 => x"0c30c3",
   40505 => x"0c30c3",
   40506 => x"0c30c3",
   40507 => x"0c30c3",
   40508 => x"0c30c3",
   40509 => x"0c30c3",
   40510 => x"0c30c3",
   40511 => x"0c30c3",
   40512 => x"0c30c3",
   40513 => x"0c30c3",
   40514 => x"0c30c3",
   40515 => x"0c30c3",
   40516 => x"0c30c3",
   40517 => x"0c30c3",
   40518 => x"0c30c3",
   40519 => x"0c30c3",
   40520 => x"0c30c3",
   40521 => x"0c30c3",
   40522 => x"0c30c3",
   40523 => x"0c30c3",
   40524 => x"0c30c3",
   40525 => x"0c30c3",
   40526 => x"0c30c3",
   40527 => x"0c30c3",
   40528 => x"0c30c3",
   40529 => x"0c30c3",
   40530 => x"0c30c3",
   40531 => x"0d7aea",
   40532 => x"aaaaaa",
   40533 => x"aaaaaa",
   40534 => x"aaaaaa",
   40535 => x"ffffff",
   40536 => x"ffffff",
   40537 => x"ffffff",
   40538 => x"ffffff",
   40539 => x"ffffff",
   40540 => x"ffffff",
   40541 => x"ffffff",
   40542 => x"ffffff",
   40543 => x"ffffff",
   40544 => x"ffffff",
   40545 => x"ffffff",
   40546 => x"ffffff",
   40547 => x"ffffff",
   40548 => x"ffffff",
   40549 => x"fffa95",
   40550 => x"abffff",
   40551 => x"ffffff",
   40552 => x"ffffff",
   40553 => x"ffffff",
   40554 => x"ffffff",
   40555 => x"ffffff",
   40556 => x"ffffff",
   40557 => x"ffffff",
   40558 => x"ffffff",
   40559 => x"ffffff",
   40560 => x"ffffff",
   40561 => x"fffb8c",
   40562 => x"30c30c",
   40563 => x"30c30c",
   40564 => x"30c30c",
   40565 => x"30c30c",
   40566 => x"30c30c",
   40567 => x"30c30c",
   40568 => x"30c30c",
   40569 => x"30c30c",
   40570 => x"30c30c",
   40571 => x"30c30c",
   40572 => x"30c30c",
   40573 => x"208208",
   40574 => x"208208",
   40575 => x"208208",
   40576 => x"208208",
   40577 => x"208208",
   40578 => x"208208",
   40579 => x"208208",
   40580 => x"208208",
   40581 => x"208208",
   40582 => x"208208",
   40583 => x"208208",
   40584 => x"208208",
   40585 => x"208208",
   40586 => x"208208",
   40587 => x"208208",
   40588 => x"208208",
   40589 => x"208208",
   40590 => x"208208",
   40591 => x"208208",
   40592 => x"208208",
   40593 => x"208208",
   40594 => x"208208",
   40595 => x"208104",
   40596 => x"104104",
   40597 => x"104104",
   40598 => x"104104",
   40599 => x"104104",
   40600 => x"104104",
   40601 => x"104104",
   40602 => x"104104",
   40603 => x"104104",
   40604 => x"104104",
   40605 => x"104104",
   40606 => x"104104",
   40607 => x"104104",
   40608 => x"104104",
   40609 => x"104104",
   40610 => x"104104",
   40611 => x"104104",
   40612 => x"104104",
   40613 => x"104104",
   40614 => x"104104",
   40615 => x"104104",
   40616 => x"104104",
   40617 => x"104104",
   40618 => x"104000",
   40619 => x"000000",
   40620 => x"000000",
   40621 => x"000000",
   40622 => x"000000",
   40623 => x"000000",
   40624 => x"000000",
   40625 => x"000000",
   40626 => x"000000",
   40627 => x"000000",
   40628 => x"000000",
   40629 => x"00057f",
   40630 => x"ffffff",
   40631 => x"ffffff",
   40632 => x"ffffff",
   40633 => x"fffa80",
   40634 => x"00002a",
   40635 => x"ffffff",
   40636 => x"ffffff",
   40637 => x"ffffff",
   40638 => x"ffffff",
   40639 => x"000000",
   40640 => x"ffffff",
   40641 => x"ffffff",
   40642 => x"ffffff",
   40643 => x"ffffff",
   40644 => x"ffffff",
   40645 => x"ffffff",
   40646 => x"ffffff",
   40647 => x"ffffff",
   40648 => x"ffffff",
   40649 => x"ffffff",
   40650 => x"ffffff",
   40651 => x"ffffff",
   40652 => x"ffffff",
   40653 => x"ffffff",
   40654 => x"ffffff",
   40655 => x"ffffff",
   40656 => x"ffffff",
   40657 => x"fd70c3",
   40658 => x"0c30c3",
   40659 => x"0c30c3",
   40660 => x"0c30c3",
   40661 => x"0c30c3",
   40662 => x"0c30c3",
   40663 => x"0c30c3",
   40664 => x"0c30c3",
   40665 => x"0c30c3",
   40666 => x"0c30c3",
   40667 => x"0c30c3",
   40668 => x"0c30c3",
   40669 => x"0c30c3",
   40670 => x"0c30c3",
   40671 => x"0c30c3",
   40672 => x"0c30c3",
   40673 => x"0c30c3",
   40674 => x"0c30c3",
   40675 => x"0c30c3",
   40676 => x"0c30c3",
   40677 => x"0c30c3",
   40678 => x"0c30c3",
   40679 => x"0c30c3",
   40680 => x"0c30c3",
   40681 => x"0c30c3",
   40682 => x"0c30c3",
   40683 => x"0c30c3",
   40684 => x"0c30c3",
   40685 => x"0c30c3",
   40686 => x"0c30c3",
   40687 => x"0c30c3",
   40688 => x"0c30c3",
   40689 => x"0c30c3",
   40690 => x"0c30c3",
   40691 => x"5ebfd5",
   40692 => x"555555",
   40693 => x"555555",
   40694 => x"555555",
   40695 => x"56aabf",
   40696 => x"ffffff",
   40697 => x"ffffff",
   40698 => x"ffffff",
   40699 => x"ffffff",
   40700 => x"ffffff",
   40701 => x"ffffff",
   40702 => x"ffffff",
   40703 => x"ffffff",
   40704 => x"ffffff",
   40705 => x"ffffff",
   40706 => x"ffffff",
   40707 => x"ffffff",
   40708 => x"ffffff",
   40709 => x"fffa95",
   40710 => x"abffff",
   40711 => x"ffffff",
   40712 => x"ffffff",
   40713 => x"ffffff",
   40714 => x"ffffff",
   40715 => x"ffffff",
   40716 => x"ffffff",
   40717 => x"ffffff",
   40718 => x"ffffff",
   40719 => x"ffffff",
   40720 => x"ffffff",
   40721 => x"fffb8c",
   40722 => x"30c30c",
   40723 => x"30c30c",
   40724 => x"30c30c",
   40725 => x"30c30c",
   40726 => x"30c30c",
   40727 => x"30c30c",
   40728 => x"30c30c",
   40729 => x"30c30c",
   40730 => x"30c30c",
   40731 => x"30c30c",
   40732 => x"30c30c",
   40733 => x"208208",
   40734 => x"208208",
   40735 => x"208208",
   40736 => x"208208",
   40737 => x"208208",
   40738 => x"208208",
   40739 => x"208208",
   40740 => x"208208",
   40741 => x"208208",
   40742 => x"208208",
   40743 => x"208208",
   40744 => x"208208",
   40745 => x"208208",
   40746 => x"208208",
   40747 => x"208208",
   40748 => x"208208",
   40749 => x"208208",
   40750 => x"208208",
   40751 => x"208208",
   40752 => x"208208",
   40753 => x"208208",
   40754 => x"208208",
   40755 => x"208104",
   40756 => x"104104",
   40757 => x"104104",
   40758 => x"104104",
   40759 => x"104104",
   40760 => x"104104",
   40761 => x"104104",
   40762 => x"104104",
   40763 => x"104104",
   40764 => x"104104",
   40765 => x"104104",
   40766 => x"104104",
   40767 => x"104104",
   40768 => x"104104",
   40769 => x"104104",
   40770 => x"104104",
   40771 => x"104104",
   40772 => x"104104",
   40773 => x"104104",
   40774 => x"104104",
   40775 => x"104104",
   40776 => x"104104",
   40777 => x"104104",
   40778 => x"104000",
   40779 => x"000000",
   40780 => x"000000",
   40781 => x"000000",
   40782 => x"000000",
   40783 => x"000000",
   40784 => x"000000",
   40785 => x"000000",
   40786 => x"000000",
   40787 => x"000000",
   40788 => x"000000",
   40789 => x"00057f",
   40790 => x"ffffff",
   40791 => x"ffffff",
   40792 => x"ffffff",
   40793 => x"ffffd5",
   40794 => x"000015",
   40795 => x"ffffff",
   40796 => x"ffffff",
   40797 => x"ffffff",
   40798 => x"ffffff",
   40799 => x"000000",
   40800 => x"ffffff",
   40801 => x"ffffff",
   40802 => x"ffffff",
   40803 => x"ffffff",
   40804 => x"ffffff",
   40805 => x"ffffff",
   40806 => x"ffffff",
   40807 => x"ffffff",
   40808 => x"ffffff",
   40809 => x"ffffff",
   40810 => x"ffffff",
   40811 => x"ffffff",
   40812 => x"ffffff",
   40813 => x"ffffff",
   40814 => x"ffffff",
   40815 => x"ffffff",
   40816 => x"ffffff",
   40817 => x"fff5c3",
   40818 => x"0c30c3",
   40819 => x"0c30c3",
   40820 => x"0c30c3",
   40821 => x"0c30c3",
   40822 => x"0c30c3",
   40823 => x"0c30c3",
   40824 => x"0c30c3",
   40825 => x"0c30c3",
   40826 => x"0c30c3",
   40827 => x"0c30c3",
   40828 => x"0c30c3",
   40829 => x"0c30c3",
   40830 => x"0c30c3",
   40831 => x"0c30c3",
   40832 => x"0c30c3",
   40833 => x"0c30c3",
   40834 => x"0c30c3",
   40835 => x"0c30c3",
   40836 => x"0c30c3",
   40837 => x"0c30c3",
   40838 => x"0c30c3",
   40839 => x"0c30c3",
   40840 => x"0c30c3",
   40841 => x"0c30c3",
   40842 => x"0c30c3",
   40843 => x"0c30c3",
   40844 => x"0c30c3",
   40845 => x"0c30c3",
   40846 => x"0c30c3",
   40847 => x"0c30c3",
   40848 => x"0c30c3",
   40849 => x"0c30c3",
   40850 => x"0c30c3",
   40851 => x"affa80",
   40852 => x"000000",
   40853 => x"000000",
   40854 => x"000000",
   40855 => x"000015",
   40856 => x"abffff",
   40857 => x"ffffff",
   40858 => x"ffffff",
   40859 => x"ffffff",
   40860 => x"ffffff",
   40861 => x"ffffff",
   40862 => x"ffffff",
   40863 => x"ffffff",
   40864 => x"ffffff",
   40865 => x"ffffff",
   40866 => x"ffffff",
   40867 => x"ffffff",
   40868 => x"ffffff",
   40869 => x"fffa95",
   40870 => x"abffff",
   40871 => x"ffffff",
   40872 => x"ffffff",
   40873 => x"ffffff",
   40874 => x"ffffff",
   40875 => x"ffffff",
   40876 => x"ffffff",
   40877 => x"ffffff",
   40878 => x"ffffff",
   40879 => x"ffffff",
   40880 => x"ffffff",
   40881 => x"fffb8c",
   40882 => x"30c30c",
   40883 => x"30c30c",
   40884 => x"30c30c",
   40885 => x"30c30c",
   40886 => x"30c30c",
   40887 => x"30c30c",
   40888 => x"30c30c",
   40889 => x"30c30c",
   40890 => x"30c30c",
   40891 => x"30c30c",
   40892 => x"30c30c",
   40893 => x"208208",
   40894 => x"208208",
   40895 => x"208208",
   40896 => x"208208",
   40897 => x"208208",
   40898 => x"208208",
   40899 => x"208208",
   40900 => x"208208",
   40901 => x"208208",
   40902 => x"208208",
   40903 => x"208208",
   40904 => x"208208",
   40905 => x"208208",
   40906 => x"208208",
   40907 => x"208208",
   40908 => x"208208",
   40909 => x"208208",
   40910 => x"208208",
   40911 => x"208208",
   40912 => x"208208",
   40913 => x"208208",
   40914 => x"208208",
   40915 => x"208104",
   40916 => x"104104",
   40917 => x"104104",
   40918 => x"104104",
   40919 => x"104104",
   40920 => x"104104",
   40921 => x"104104",
   40922 => x"104104",
   40923 => x"104104",
   40924 => x"104104",
   40925 => x"104104",
   40926 => x"104104",
   40927 => x"104104",
   40928 => x"104104",
   40929 => x"104104",
   40930 => x"104104",
   40931 => x"104104",
   40932 => x"104104",
   40933 => x"104104",
   40934 => x"104104",
   40935 => x"104104",
   40936 => x"104104",
   40937 => x"104104",
   40938 => x"104000",
   40939 => x"000000",
   40940 => x"000000",
   40941 => x"000000",
   40942 => x"000000",
   40943 => x"000000",
   40944 => x"000000",
   40945 => x"000000",
   40946 => x"000000",
   40947 => x"000000",
   40948 => x"000000",
   40949 => x"00057f",
   40950 => x"ffffff",
   40951 => x"ffffff",
   40952 => x"ffffff",
   40953 => x"ffffea",
   40954 => x"000000",
   40955 => x"abffff",
   40956 => x"ffffff",
   40957 => x"ffffff",
   40958 => x"ffffff",
   40959 => x"000000",
   40960 => x"ffffff",
   40961 => x"ffffff",
   40962 => x"ffffff",
   40963 => x"ffffff",
   40964 => x"ffffff",
   40965 => x"ffffff",
   40966 => x"ffffff",
   40967 => x"ffffff",
   40968 => x"ffffff",
   40969 => x"ffffff",
   40970 => x"ffffff",
   40971 => x"ffffff",
   40972 => x"ffffff",
   40973 => x"ffffff",
   40974 => x"ffffff",
   40975 => x"ffffff",
   40976 => x"ffffff",
   40977 => x"ffffd7",
   40978 => x"0c30c3",
   40979 => x"0c30c3",
   40980 => x"0c30c3",
   40981 => x"0c30c3",
   40982 => x"0c30c3",
   40983 => x"0c30c3",
   40984 => x"0c30c3",
   40985 => x"0c30c3",
   40986 => x"0c30c3",
   40987 => x"0c30c3",
   40988 => x"0c30c3",
   40989 => x"0c30c3",
   40990 => x"0c30c3",
   40991 => x"0c30c3",
   40992 => x"0c30c3",
   40993 => x"0c30c3",
   40994 => x"0c30c3",
   40995 => x"0c30c3",
   40996 => x"0c30c3",
   40997 => x"0c30c3",
   40998 => x"0c30c3",
   40999 => x"0c30c3",
   41000 => x"0c30c3",
   41001 => x"0c30c3",
   41002 => x"0c30c3",
   41003 => x"0c30c3",
   41004 => x"0c30c3",
   41005 => x"0c30c3",
   41006 => x"0c30c3",
   41007 => x"0c30c3",
   41008 => x"0c30c3",
   41009 => x"0c30c3",
   41010 => x"0c30eb",
   41011 => x"fffa80",
   41012 => x"000000",
   41013 => x"000000",
   41014 => x"000000",
   41015 => x"000000",
   41016 => x"56afff",
   41017 => x"ffffff",
   41018 => x"ffffff",
   41019 => x"ffffff",
   41020 => x"ffffff",
   41021 => x"ffffff",
   41022 => x"ffffff",
   41023 => x"ffffff",
   41024 => x"ffffff",
   41025 => x"ffffff",
   41026 => x"ffffff",
   41027 => x"ffffff",
   41028 => x"ffffff",
   41029 => x"fffa95",
   41030 => x"abffff",
   41031 => x"ffffff",
   41032 => x"ffffff",
   41033 => x"ffffff",
   41034 => x"ffffff",
   41035 => x"ffffff",
   41036 => x"ffffff",
   41037 => x"ffffff",
   41038 => x"ffffff",
   41039 => x"ffffff",
   41040 => x"ffffff",
   41041 => x"fffb8c",
   41042 => x"30c30c",
   41043 => x"30c30c",
   41044 => x"30c30c",
   41045 => x"30c30c",
   41046 => x"30c30c",
   41047 => x"30c30c",
   41048 => x"30c30c",
   41049 => x"30c30c",
   41050 => x"30c30c",
   41051 => x"30c30c",
   41052 => x"30c30c",
   41053 => x"208208",
   41054 => x"208208",
   41055 => x"208208",
   41056 => x"208208",
   41057 => x"208208",
   41058 => x"208208",
   41059 => x"208208",
   41060 => x"208208",
   41061 => x"208208",
   41062 => x"208208",
   41063 => x"208208",
   41064 => x"208208",
   41065 => x"208208",
   41066 => x"208208",
   41067 => x"208208",
   41068 => x"208208",
   41069 => x"208208",
   41070 => x"208208",
   41071 => x"208208",
   41072 => x"208208",
   41073 => x"208208",
   41074 => x"208208",
   41075 => x"208104",
   41076 => x"104104",
   41077 => x"104104",
   41078 => x"104104",
   41079 => x"104104",
   41080 => x"104104",
   41081 => x"104104",
   41082 => x"104104",
   41083 => x"104104",
   41084 => x"104104",
   41085 => x"104104",
   41086 => x"104104",
   41087 => x"104104",
   41088 => x"104104",
   41089 => x"104104",
   41090 => x"104104",
   41091 => x"104104",
   41092 => x"104104",
   41093 => x"104104",
   41094 => x"104104",
   41095 => x"104104",
   41096 => x"104104",
   41097 => x"104104",
   41098 => x"104000",
   41099 => x"000000",
   41100 => x"000000",
   41101 => x"000000",
   41102 => x"000000",
   41103 => x"000000",
   41104 => x"000000",
   41105 => x"000000",
   41106 => x"000000",
   41107 => x"000000",
   41108 => x"000000",
   41109 => x"00057f",
   41110 => x"ffffff",
   41111 => x"ffffff",
   41112 => x"ffffff",
   41113 => x"ffffff",
   41114 => x"540000",
   41115 => x"02afff",
   41116 => x"ffffff",
   41117 => x"ffffff",
   41118 => x"ffffea",
   41119 => x"000000",
   41120 => x"ffffff",
   41121 => x"ffffff",
   41122 => x"ffffff",
   41123 => x"ffffff",
   41124 => x"ffffff",
   41125 => x"ffffff",
   41126 => x"ffffff",
   41127 => x"ffffff",
   41128 => x"ffffff",
   41129 => x"ffffff",
   41130 => x"ffffff",
   41131 => x"ffffff",
   41132 => x"ffffff",
   41133 => x"ffffff",
   41134 => x"ffffff",
   41135 => x"ffffff",
   41136 => x"ffffff",
   41137 => x"ffffff",
   41138 => x"5c30c3",
   41139 => x"0c30c3",
   41140 => x"0c30c3",
   41141 => x"0c30c3",
   41142 => x"0c30c3",
   41143 => x"0c30c3",
   41144 => x"0c30c3",
   41145 => x"0c30c3",
   41146 => x"0c30c3",
   41147 => x"0c30c3",
   41148 => x"0c30c3",
   41149 => x"0c30c3",
   41150 => x"0c30c3",
   41151 => x"0c30c3",
   41152 => x"0c30c3",
   41153 => x"0c30c3",
   41154 => x"0c30c3",
   41155 => x"0c30c3",
   41156 => x"0c30c3",
   41157 => x"0c30c3",
   41158 => x"0c30c3",
   41159 => x"0c30c3",
   41160 => x"0c30c3",
   41161 => x"0c30c3",
   41162 => x"0c30c3",
   41163 => x"0c30c3",
   41164 => x"0c30c3",
   41165 => x"0c30c3",
   41166 => x"0c30c3",
   41167 => x"0c30c3",
   41168 => x"0c30c3",
   41169 => x"0c30c3",
   41170 => x"0c3aff",
   41171 => x"fffa80",
   41172 => x"000015",
   41173 => x"aaaaaa",
   41174 => x"aaa555",
   41175 => x"540000",
   41176 => x"015abf",
   41177 => x"ffffff",
   41178 => x"ffffff",
   41179 => x"ffffff",
   41180 => x"ffffff",
   41181 => x"ffffff",
   41182 => x"ffffff",
   41183 => x"ffffff",
   41184 => x"ffffff",
   41185 => x"ffffff",
   41186 => x"ffffff",
   41187 => x"ffffff",
   41188 => x"ffffff",
   41189 => x"fffa95",
   41190 => x"abffff",
   41191 => x"ffffff",
   41192 => x"ffffff",
   41193 => x"ffffff",
   41194 => x"ffffff",
   41195 => x"ffffff",
   41196 => x"ffffff",
   41197 => x"ffffff",
   41198 => x"ffffff",
   41199 => x"ffffff",
   41200 => x"ffffff",
   41201 => x"fffb8c",
   41202 => x"30c30c",
   41203 => x"30c30c",
   41204 => x"30c30c",
   41205 => x"30c30c",
   41206 => x"30c30c",
   41207 => x"30c30c",
   41208 => x"30c30c",
   41209 => x"30c30c",
   41210 => x"30c30c",
   41211 => x"30c30c",
   41212 => x"30c30c",
   41213 => x"208208",
   41214 => x"208208",
   41215 => x"208208",
   41216 => x"208208",
   41217 => x"208208",
   41218 => x"208208",
   41219 => x"208208",
   41220 => x"208208",
   41221 => x"208208",
   41222 => x"208208",
   41223 => x"208208",
   41224 => x"208208",
   41225 => x"208208",
   41226 => x"208208",
   41227 => x"208208",
   41228 => x"208208",
   41229 => x"208208",
   41230 => x"208208",
   41231 => x"208208",
   41232 => x"208208",
   41233 => x"208208",
   41234 => x"208208",
   41235 => x"208104",
   41236 => x"104104",
   41237 => x"104104",
   41238 => x"104104",
   41239 => x"104104",
   41240 => x"104104",
   41241 => x"104104",
   41242 => x"104104",
   41243 => x"104104",
   41244 => x"104104",
   41245 => x"104104",
   41246 => x"104104",
   41247 => x"104104",
   41248 => x"104104",
   41249 => x"104104",
   41250 => x"104104",
   41251 => x"104104",
   41252 => x"104104",
   41253 => x"104104",
   41254 => x"104104",
   41255 => x"104104",
   41256 => x"104104",
   41257 => x"104104",
   41258 => x"104000",
   41259 => x"000000",
   41260 => x"000000",
   41261 => x"000000",
   41262 => x"000000",
   41263 => x"000000",
   41264 => x"000000",
   41265 => x"000000",
   41266 => x"000000",
   41267 => x"000000",
   41268 => x"000000",
   41269 => x"00057f",
   41270 => x"ffffff",
   41271 => x"ffffff",
   41272 => x"ffffff",
   41273 => x"ffffff",
   41274 => x"a95000",
   41275 => x"00056a",
   41276 => x"ffffff",
   41277 => x"ffffff",
   41278 => x"fffaaa",
   41279 => x"000000",
   41280 => x"ffffff",
   41281 => x"ffffff",
   41282 => x"ffffff",
   41283 => x"ffffff",
   41284 => x"ffffff",
   41285 => x"ffffff",
   41286 => x"ffffff",
   41287 => x"ffffff",
   41288 => x"ffffff",
   41289 => x"ffffff",
   41290 => x"ffffff",
   41291 => x"ffffff",
   41292 => x"ffffff",
   41293 => x"ffffff",
   41294 => x"ffffff",
   41295 => x"ffffff",
   41296 => x"ffffff",
   41297 => x"ffffff",
   41298 => x"fd70c3",
   41299 => x"0c30c3",
   41300 => x"0c30c3",
   41301 => x"0c30c3",
   41302 => x"0c30c3",
   41303 => x"0c30c3",
   41304 => x"0c30c3",
   41305 => x"0c30c3",
   41306 => x"0c30c3",
   41307 => x"0c30c3",
   41308 => x"0c30c3",
   41309 => x"0c30c3",
   41310 => x"0c30c3",
   41311 => x"0c30c3",
   41312 => x"0c30c3",
   41313 => x"0c30c3",
   41314 => x"0c30c3",
   41315 => x"0c30c3",
   41316 => x"0c30c3",
   41317 => x"0c30c3",
   41318 => x"0c30c3",
   41319 => x"0c30c3",
   41320 => x"0c30c3",
   41321 => x"0c30c3",
   41322 => x"0c30c3",
   41323 => x"0c30c3",
   41324 => x"0c30c3",
   41325 => x"0c30c3",
   41326 => x"0c30c3",
   41327 => x"0c30c3",
   41328 => x"0c30c3",
   41329 => x"0c30c3",
   41330 => x"0ebfff",
   41331 => x"fffa80",
   41332 => x"00003f",
   41333 => x"ffffff",
   41334 => x"ffffff",
   41335 => x"fd5000",
   41336 => x"00057f",
   41337 => x"ffffff",
   41338 => x"ffffff",
   41339 => x"ffffff",
   41340 => x"ffffff",
   41341 => x"ffffff",
   41342 => x"ffffff",
   41343 => x"ffffff",
   41344 => x"ffffff",
   41345 => x"ffffff",
   41346 => x"ffffff",
   41347 => x"ffffff",
   41348 => x"ffffff",
   41349 => x"fffa95",
   41350 => x"abffff",
   41351 => x"ffffff",
   41352 => x"ffffff",
   41353 => x"ffffff",
   41354 => x"ffffff",
   41355 => x"ffffff",
   41356 => x"ffffff",
   41357 => x"ffffff",
   41358 => x"ffffff",
   41359 => x"ffffff",
   41360 => x"ffffff",
   41361 => x"fffb8c",
   41362 => x"30c30c",
   41363 => x"30c30c",
   41364 => x"30c30c",
   41365 => x"30c30c",
   41366 => x"30c30c",
   41367 => x"30c30c",
   41368 => x"30c30c",
   41369 => x"30c30c",
   41370 => x"30c30c",
   41371 => x"30c30c",
   41372 => x"30c30c",
   41373 => x"208208",
   41374 => x"208208",
   41375 => x"208208",
   41376 => x"208208",
   41377 => x"208208",
   41378 => x"208208",
   41379 => x"208208",
   41380 => x"208208",
   41381 => x"208208",
   41382 => x"208208",
   41383 => x"208208",
   41384 => x"208208",
   41385 => x"208208",
   41386 => x"208208",
   41387 => x"208208",
   41388 => x"208208",
   41389 => x"208208",
   41390 => x"208208",
   41391 => x"208208",
   41392 => x"208208",
   41393 => x"208208",
   41394 => x"208208",
   41395 => x"208104",
   41396 => x"104104",
   41397 => x"104104",
   41398 => x"104104",
   41399 => x"104104",
   41400 => x"104104",
   41401 => x"104104",
   41402 => x"104104",
   41403 => x"104104",
   41404 => x"104104",
   41405 => x"104104",
   41406 => x"104104",
   41407 => x"104104",
   41408 => x"104104",
   41409 => x"104104",
   41410 => x"104104",
   41411 => x"104104",
   41412 => x"104104",
   41413 => x"104104",
   41414 => x"104104",
   41415 => x"104104",
   41416 => x"104104",
   41417 => x"104104",
   41418 => x"104000",
   41419 => x"000000",
   41420 => x"000000",
   41421 => x"000000",
   41422 => x"000000",
   41423 => x"000000",
   41424 => x"000000",
   41425 => x"000000",
   41426 => x"000000",
   41427 => x"000000",
   41428 => x"000000",
   41429 => x"00057f",
   41430 => x"ffffff",
   41431 => x"ffffff",
   41432 => x"ffffff",
   41433 => x"ffffff",
   41434 => x"fea540",
   41435 => x"000000",
   41436 => x"56aaaa",
   41437 => x"feaaaa",
   41438 => x"a95000",
   41439 => x"000000",
   41440 => x"ffffff",
   41441 => x"ffffff",
   41442 => x"ffffff",
   41443 => x"ffffff",
   41444 => x"ffffff",
   41445 => x"ffffff",
   41446 => x"ffffff",
   41447 => x"ffffff",
   41448 => x"ffffff",
   41449 => x"ffffff",
   41450 => x"ffffff",
   41451 => x"ffffff",
   41452 => x"ffffff",
   41453 => x"ffffff",
   41454 => x"ffffff",
   41455 => x"ffffff",
   41456 => x"ffffff",
   41457 => x"ffffff",
   41458 => x"fff5c3",
   41459 => x"0c30c3",
   41460 => x"0c30c3",
   41461 => x"0c30c3",
   41462 => x"0c30c3",
   41463 => x"0c30c3",
   41464 => x"0c30c3",
   41465 => x"0c30c3",
   41466 => x"0c30c3",
   41467 => x"0c30c3",
   41468 => x"0c30c3",
   41469 => x"0c30c3",
   41470 => x"0c30c3",
   41471 => x"0c30c3",
   41472 => x"0c30c3",
   41473 => x"0c30c3",
   41474 => x"0c30c3",
   41475 => x"0c30c3",
   41476 => x"0c30c3",
   41477 => x"0c30c3",
   41478 => x"0c30c3",
   41479 => x"0c30c3",
   41480 => x"0c30c3",
   41481 => x"0c30c3",
   41482 => x"0c30c3",
   41483 => x"0c30c3",
   41484 => x"0c30c3",
   41485 => x"0c30c3",
   41486 => x"0c30c3",
   41487 => x"0c30c3",
   41488 => x"0c30c3",
   41489 => x"0c30d7",
   41490 => x"afffff",
   41491 => x"fffa80",
   41492 => x"00003f",
   41493 => x"ffffff",
   41494 => x"ffffff",
   41495 => x"fff540",
   41496 => x"00056a",
   41497 => x"ffffff",
   41498 => x"ffffff",
   41499 => x"ffffff",
   41500 => x"ffffff",
   41501 => x"ffffff",
   41502 => x"ffffff",
   41503 => x"ffffff",
   41504 => x"ffffff",
   41505 => x"ffffff",
   41506 => x"ffffff",
   41507 => x"ffffff",
   41508 => x"ffffff",
   41509 => x"fffa95",
   41510 => x"abffff",
   41511 => x"ffffff",
   41512 => x"ffffff",
   41513 => x"ffffff",
   41514 => x"ffffff",
   41515 => x"ffffff",
   41516 => x"ffffff",
   41517 => x"ffffff",
   41518 => x"ffffff",
   41519 => x"ffffff",
   41520 => x"ffffff",
   41521 => x"fffb8c",
   41522 => x"30c30c",
   41523 => x"30c30c",
   41524 => x"30c30c",
   41525 => x"30c30c",
   41526 => x"30c30c",
   41527 => x"30c30c",
   41528 => x"30c30c",
   41529 => x"30c30c",
   41530 => x"30c30c",
   41531 => x"30c30c",
   41532 => x"30c30c",
   41533 => x"208208",
   41534 => x"208208",
   41535 => x"208208",
   41536 => x"208208",
   41537 => x"208208",
   41538 => x"208208",
   41539 => x"208208",
   41540 => x"208208",
   41541 => x"208208",
   41542 => x"208208",
   41543 => x"208208",
   41544 => x"208208",
   41545 => x"208208",
   41546 => x"208208",
   41547 => x"208208",
   41548 => x"208208",
   41549 => x"208208",
   41550 => x"208208",
   41551 => x"208208",
   41552 => x"208208",
   41553 => x"208208",
   41554 => x"208208",
   41555 => x"208104",
   41556 => x"104104",
   41557 => x"104104",
   41558 => x"104104",
   41559 => x"104104",
   41560 => x"104104",
   41561 => x"104104",
   41562 => x"104104",
   41563 => x"104104",
   41564 => x"104104",
   41565 => x"104104",
   41566 => x"104104",
   41567 => x"104104",
   41568 => x"104104",
   41569 => x"104104",
   41570 => x"104104",
   41571 => x"104104",
   41572 => x"104104",
   41573 => x"104104",
   41574 => x"104104",
   41575 => x"104104",
   41576 => x"104104",
   41577 => x"104104",
   41578 => x"104000",
   41579 => x"000000",
   41580 => x"000000",
   41581 => x"000000",
   41582 => x"000000",
   41583 => x"000000",
   41584 => x"000000",
   41585 => x"000000",
   41586 => x"000000",
   41587 => x"000000",
   41588 => x"000000",
   41589 => x"00057f",
   41590 => x"ffffff",
   41591 => x"ffffff",
   41592 => x"ffffff",
   41593 => x"ffffff",
   41594 => x"fffa95",
   41595 => x"000000",
   41596 => x"000000",
   41597 => x"000000",
   41598 => x"000000",
   41599 => x"00056a",
   41600 => x"ffffff",
   41601 => x"ffffff",
   41602 => x"ffffff",
   41603 => x"ffffff",
   41604 => x"ffffff",
   41605 => x"ffffff",
   41606 => x"ffffff",
   41607 => x"ffffff",
   41608 => x"ffffff",
   41609 => x"ffffff",
   41610 => x"ffffff",
   41611 => x"ffffff",
   41612 => x"ffffff",
   41613 => x"ffffff",
   41614 => x"ffffff",
   41615 => x"ffffff",
   41616 => x"ffffff",
   41617 => x"ffffff",
   41618 => x"ffffeb",
   41619 => x"0c30c3",
   41620 => x"0c30c3",
   41621 => x"0c30c3",
   41622 => x"0c30c3",
   41623 => x"0c30c3",
   41624 => x"0c30c3",
   41625 => x"0c30c3",
   41626 => x"0c30c3",
   41627 => x"0c30c3",
   41628 => x"0c30c3",
   41629 => x"0c30c3",
   41630 => x"0c30c3",
   41631 => x"0c30c3",
   41632 => x"0c30c3",
   41633 => x"0c30c3",
   41634 => x"0c30c3",
   41635 => x"0c30c3",
   41636 => x"0c30c3",
   41637 => x"0c30c3",
   41638 => x"0c30c3",
   41639 => x"0c30c3",
   41640 => x"0c30c3",
   41641 => x"0c30c3",
   41642 => x"0c30c3",
   41643 => x"0c30c3",
   41644 => x"0c30c3",
   41645 => x"0c30c3",
   41646 => x"0c30c3",
   41647 => x"0c30c3",
   41648 => x"0c30c3",
   41649 => x"0c35eb",
   41650 => x"ffffff",
   41651 => x"fffa80",
   41652 => x"00003f",
   41653 => x"ffffff",
   41654 => x"ffffff",
   41655 => x"fffa80",
   41656 => x"00056a",
   41657 => x"ffffff",
   41658 => x"ffffff",
   41659 => x"ffffff",
   41660 => x"ffffff",
   41661 => x"ffffff",
   41662 => x"ffffff",
   41663 => x"ffffff",
   41664 => x"ffffff",
   41665 => x"ffffff",
   41666 => x"ffffff",
   41667 => x"ffffff",
   41668 => x"ffffff",
   41669 => x"fffa95",
   41670 => x"abffff",
   41671 => x"ffffff",
   41672 => x"ffffff",
   41673 => x"ffffff",
   41674 => x"ffffff",
   41675 => x"ffffff",
   41676 => x"ffffff",
   41677 => x"ffffff",
   41678 => x"ffffff",
   41679 => x"ffffff",
   41680 => x"ffffff",
   41681 => x"fffb8c",
   41682 => x"30c30c",
   41683 => x"30c30c",
   41684 => x"30c30c",
   41685 => x"30c30c",
   41686 => x"30c30c",
   41687 => x"30c30c",
   41688 => x"30c30c",
   41689 => x"30c30c",
   41690 => x"30c30c",
   41691 => x"30c30c",
   41692 => x"30c30c",
   41693 => x"208208",
   41694 => x"208208",
   41695 => x"208208",
   41696 => x"208208",
   41697 => x"208208",
   41698 => x"208208",
   41699 => x"208208",
   41700 => x"208208",
   41701 => x"208208",
   41702 => x"208208",
   41703 => x"208208",
   41704 => x"208208",
   41705 => x"208208",
   41706 => x"208208",
   41707 => x"208208",
   41708 => x"208208",
   41709 => x"208208",
   41710 => x"208208",
   41711 => x"208208",
   41712 => x"208208",
   41713 => x"208208",
   41714 => x"208208",
   41715 => x"208104",
   41716 => x"104104",
   41717 => x"104104",
   41718 => x"104104",
   41719 => x"104104",
   41720 => x"104104",
   41721 => x"104104",
   41722 => x"104104",
   41723 => x"104104",
   41724 => x"104104",
   41725 => x"104104",
   41726 => x"104104",
   41727 => x"104104",
   41728 => x"104104",
   41729 => x"104104",
   41730 => x"104104",
   41731 => x"104104",
   41732 => x"104104",
   41733 => x"104104",
   41734 => x"104104",
   41735 => x"104104",
   41736 => x"104104",
   41737 => x"104104",
   41738 => x"104000",
   41739 => x"000000",
   41740 => x"000000",
   41741 => x"000000",
   41742 => x"000000",
   41743 => x"000000",
   41744 => x"000000",
   41745 => x"000000",
   41746 => x"000000",
   41747 => x"000000",
   41748 => x"000000",
   41749 => x"00057f",
   41750 => x"ffffff",
   41751 => x"ffffff",
   41752 => x"ffffff",
   41753 => x"ffffff",
   41754 => x"ffffff",
   41755 => x"a95000",
   41756 => x"000000",
   41757 => x"000000",
   41758 => x"000000",
   41759 => x"56afff",
   41760 => x"ffffff",
   41761 => x"ffffff",
   41762 => x"ffffff",
   41763 => x"ffffff",
   41764 => x"ffffff",
   41765 => x"ffffff",
   41766 => x"ffffff",
   41767 => x"ffffff",
   41768 => x"ffffff",
   41769 => x"ffffff",
   41770 => x"ffffff",
   41771 => x"ffffff",
   41772 => x"ffffff",
   41773 => x"ffffff",
   41774 => x"ffffff",
   41775 => x"ffffff",
   41776 => x"ffffff",
   41777 => x"ffffff",
   41778 => x"ffffff",
   41779 => x"ac30c3",
   41780 => x"0c30c3",
   41781 => x"0c30c3",
   41782 => x"0c30c3",
   41783 => x"0c30c3",
   41784 => x"0c30c3",
   41785 => x"0c30c3",
   41786 => x"0c30c3",
   41787 => x"0c30c3",
   41788 => x"0c30c3",
   41789 => x"0c30c3",
   41790 => x"0c30c3",
   41791 => x"0c30c3",
   41792 => x"0c30c3",
   41793 => x"0c30c3",
   41794 => x"0c30c3",
   41795 => x"0c30c3",
   41796 => x"0c30c3",
   41797 => x"0c30c3",
   41798 => x"0c30c3",
   41799 => x"0c30c3",
   41800 => x"0c30c3",
   41801 => x"0c30c3",
   41802 => x"0c30c3",
   41803 => x"0c30c3",
   41804 => x"0c30c3",
   41805 => x"0c30c3",
   41806 => x"0c30c3",
   41807 => x"0c30c3",
   41808 => x"0c30c3",
   41809 => x"0d7aff",
   41810 => x"ffffff",
   41811 => x"fffa80",
   41812 => x"00003f",
   41813 => x"ffffff",
   41814 => x"ffffff",
   41815 => x"fffa95",
   41816 => x"00002a",
   41817 => x"ffffff",
   41818 => x"ffffff",
   41819 => x"ffffff",
   41820 => x"ffffff",
   41821 => x"ffffff",
   41822 => x"ffffff",
   41823 => x"ffffff",
   41824 => x"ffffff",
   41825 => x"ffffff",
   41826 => x"ffffff",
   41827 => x"ffffff",
   41828 => x"ffffff",
   41829 => x"fffa95",
   41830 => x"abffff",
   41831 => x"ffffff",
   41832 => x"ffffff",
   41833 => x"ffffff",
   41834 => x"ffffff",
   41835 => x"ffffff",
   41836 => x"ffffff",
   41837 => x"ffffff",
   41838 => x"ffffff",
   41839 => x"ffffff",
   41840 => x"ffffff",
   41841 => x"fffb8c",
   41842 => x"30c30c",
   41843 => x"30c30c",
   41844 => x"30c30c",
   41845 => x"30c30c",
   41846 => x"30c30c",
   41847 => x"30c30c",
   41848 => x"30c30c",
   41849 => x"30c30c",
   41850 => x"30c30c",
   41851 => x"30c30c",
   41852 => x"30c30c",
   41853 => x"208208",
   41854 => x"208208",
   41855 => x"208208",
   41856 => x"208208",
   41857 => x"208208",
   41858 => x"208208",
   41859 => x"208208",
   41860 => x"208208",
   41861 => x"208208",
   41862 => x"208208",
   41863 => x"208208",
   41864 => x"208208",
   41865 => x"208208",
   41866 => x"208208",
   41867 => x"208208",
   41868 => x"208208",
   41869 => x"208208",
   41870 => x"208208",
   41871 => x"208208",
   41872 => x"208208",
   41873 => x"208208",
   41874 => x"208208",
   41875 => x"208104",
   41876 => x"104104",
   41877 => x"104104",
   41878 => x"104104",
   41879 => x"104104",
   41880 => x"104104",
   41881 => x"104104",
   41882 => x"104104",
   41883 => x"104104",
   41884 => x"104104",
   41885 => x"104104",
   41886 => x"104104",
   41887 => x"104104",
   41888 => x"104104",
   41889 => x"104104",
   41890 => x"104104",
   41891 => x"104104",
   41892 => x"104104",
   41893 => x"104104",
   41894 => x"104104",
   41895 => x"104104",
   41896 => x"104104",
   41897 => x"104104",
   41898 => x"104000",
   41899 => x"000000",
   41900 => x"000000",
   41901 => x"000000",
   41902 => x"000000",
   41903 => x"000000",
   41904 => x"000000",
   41905 => x"000000",
   41906 => x"000000",
   41907 => x"000000",
   41908 => x"000000",
   41909 => x"00057f",
   41910 => x"ffffff",
   41911 => x"ffffff",
   41912 => x"ffffff",
   41913 => x"ffffff",
   41914 => x"ffffff",
   41915 => x"fffa95",
   41916 => x"540000",
   41917 => x"000000",
   41918 => x"01556a",
   41919 => x"ffffff",
   41920 => x"ffffff",
   41921 => x"ffffff",
   41922 => x"ffffff",
   41923 => x"ffffff",
   41924 => x"ffffff",
   41925 => x"ffffff",
   41926 => x"ffffff",
   41927 => x"ffffff",
   41928 => x"ffffff",
   41929 => x"ffffff",
   41930 => x"ffffff",
   41931 => x"ffffff",
   41932 => x"ffffff",
   41933 => x"ffffff",
   41934 => x"ffffff",
   41935 => x"ffffff",
   41936 => x"ffffff",
   41937 => x"ffffff",
   41938 => x"ffffff",
   41939 => x"feb0c3",
   41940 => x"0c30c3",
   41941 => x"0c30c3",
   41942 => x"0c30c3",
   41943 => x"0c30c3",
   41944 => x"0c30c3",
   41945 => x"0c30c3",
   41946 => x"0c30c3",
   41947 => x"0c30c3",
   41948 => x"0c30c3",
   41949 => x"0c30c3",
   41950 => x"0c30c3",
   41951 => x"0c30c3",
   41952 => x"0c30c3",
   41953 => x"0c30c3",
   41954 => x"0c30c3",
   41955 => x"0c30c3",
   41956 => x"0c30c3",
   41957 => x"0c30c3",
   41958 => x"0c30c3",
   41959 => x"0c30c3",
   41960 => x"0c30c3",
   41961 => x"0c30c3",
   41962 => x"0c30c3",
   41963 => x"0c30c3",
   41964 => x"0c30c3",
   41965 => x"0c30c3",
   41966 => x"0c30c3",
   41967 => x"0c30c3",
   41968 => x"0c30c3",
   41969 => x"5ebfff",
   41970 => x"ffffff",
   41971 => x"fffa80",
   41972 => x"00003f",
   41973 => x"ffffff",
   41974 => x"ffffff",
   41975 => x"fffa95",
   41976 => x"00056a",
   41977 => x"ffffff",
   41978 => x"ffffff",
   41979 => x"ffffff",
   41980 => x"ffffff",
   41981 => x"ffffff",
   41982 => x"ffffff",
   41983 => x"ffffff",
   41984 => x"ffffff",
   41985 => x"ffffff",
   41986 => x"ffffff",
   41987 => x"ffffff",
   41988 => x"ffffff",
   41989 => x"fffa95",
   41990 => x"abffff",
   41991 => x"ffffff",
   41992 => x"ffffff",
   41993 => x"ffffff",
   41994 => x"ffffff",
   41995 => x"ffffff",
   41996 => x"ffffff",
   41997 => x"ffffff",
   41998 => x"ffffff",
   41999 => x"ffffff",
   42000 => x"ffffff",
   42001 => x"fffb8c",
   42002 => x"30c30c",
   42003 => x"30c30c",
   42004 => x"30c30c",
   42005 => x"30c30c",
   42006 => x"30c30c",
   42007 => x"30c30c",
   42008 => x"30c30c",
   42009 => x"30c30c",
   42010 => x"30c30c",
   42011 => x"30c30c",
   42012 => x"30c30c",
   42013 => x"208208",
   42014 => x"208208",
   42015 => x"208208",
   42016 => x"208208",
   42017 => x"208208",
   42018 => x"208208",
   42019 => x"208208",
   42020 => x"208208",
   42021 => x"208208",
   42022 => x"208208",
   42023 => x"208208",
   42024 => x"208208",
   42025 => x"208208",
   42026 => x"208208",
   42027 => x"208208",
   42028 => x"208208",
   42029 => x"208208",
   42030 => x"208208",
   42031 => x"208208",
   42032 => x"208208",
   42033 => x"208208",
   42034 => x"208208",
   42035 => x"208104",
   42036 => x"104104",
   42037 => x"104104",
   42038 => x"104104",
   42039 => x"104104",
   42040 => x"104104",
   42041 => x"104104",
   42042 => x"104104",
   42043 => x"104104",
   42044 => x"104104",
   42045 => x"104104",
   42046 => x"104104",
   42047 => x"104104",
   42048 => x"104104",
   42049 => x"104104",
   42050 => x"104104",
   42051 => x"104104",
   42052 => x"104104",
   42053 => x"104104",
   42054 => x"104104",
   42055 => x"104104",
   42056 => x"104104",
   42057 => x"104104",
   42058 => x"104000",
   42059 => x"000000",
   42060 => x"000000",
   42061 => x"000000",
   42062 => x"000000",
   42063 => x"000000",
   42064 => x"000000",
   42065 => x"000000",
   42066 => x"000000",
   42067 => x"000000",
   42068 => x"000000",
   42069 => x"00057f",
   42070 => x"ffffff",
   42071 => x"ffffff",
   42072 => x"ffffff",
   42073 => x"ffffff",
   42074 => x"ffffff",
   42075 => x"ffffff",
   42076 => x"fffaaa",
   42077 => x"aaaabf",
   42078 => x"ffffff",
   42079 => x"ffffff",
   42080 => x"ffffff",
   42081 => x"ffffff",
   42082 => x"ffffff",
   42083 => x"ffffff",
   42084 => x"ffffff",
   42085 => x"ffffff",
   42086 => x"ffffff",
   42087 => x"ffffff",
   42088 => x"ffffff",
   42089 => x"ffffff",
   42090 => x"ffffff",
   42091 => x"ffffff",
   42092 => x"ffffff",
   42093 => x"ffffff",
   42094 => x"ffffff",
   42095 => x"ffffff",
   42096 => x"ffffff",
   42097 => x"ffffff",
   42098 => x"ffffff",
   42099 => x"fffad7",
   42100 => x"0c30c3",
   42101 => x"0c30c3",
   42102 => x"0c30c3",
   42103 => x"0c30c3",
   42104 => x"0c30c3",
   42105 => x"0c30c3",
   42106 => x"0c30c3",
   42107 => x"0c30c3",
   42108 => x"0c30c3",
   42109 => x"0c30c3",
   42110 => x"0c30c3",
   42111 => x"0c30c3",
   42112 => x"0c30c3",
   42113 => x"0c30c3",
   42114 => x"0c30c3",
   42115 => x"0c30c3",
   42116 => x"0c30c3",
   42117 => x"0c30c3",
   42118 => x"0c30c3",
   42119 => x"0c30c3",
   42120 => x"0c30c3",
   42121 => x"0c30c3",
   42122 => x"0c30c3",
   42123 => x"0c30c3",
   42124 => x"0c30c3",
   42125 => x"0c30c3",
   42126 => x"0c30c3",
   42127 => x"0c30c3",
   42128 => x"0c30d7",
   42129 => x"ffffff",
   42130 => x"ffffff",
   42131 => x"fffa80",
   42132 => x"00003f",
   42133 => x"ffffff",
   42134 => x"ffffff",
   42135 => x"fffa80",
   42136 => x"00056a",
   42137 => x"ffffff",
   42138 => x"ffffff",
   42139 => x"ffffff",
   42140 => x"ffffff",
   42141 => x"ffffff",
   42142 => x"ffffff",
   42143 => x"ffffff",
   42144 => x"ffffff",
   42145 => x"ffffff",
   42146 => x"ffffff",
   42147 => x"ffffff",
   42148 => x"ffffff",
   42149 => x"fffa95",
   42150 => x"abffff",
   42151 => x"ffffff",
   42152 => x"ffffff",
   42153 => x"ffffff",
   42154 => x"ffffff",
   42155 => x"ffffff",
   42156 => x"ffffff",
   42157 => x"ffffff",
   42158 => x"ffffff",
   42159 => x"ffffff",
   42160 => x"ffffff",
   42161 => x"fffb8c",
   42162 => x"30c30c",
   42163 => x"30c30c",
   42164 => x"30c30c",
   42165 => x"30c30c",
   42166 => x"30c30c",
   42167 => x"30c30c",
   42168 => x"30c30c",
   42169 => x"30c30c",
   42170 => x"30c30c",
   42171 => x"30c30c",
   42172 => x"30c30c",
   42173 => x"208208",
   42174 => x"208208",
   42175 => x"208208",
   42176 => x"208208",
   42177 => x"208208",
   42178 => x"208208",
   42179 => x"208208",
   42180 => x"208208",
   42181 => x"208208",
   42182 => x"208208",
   42183 => x"208208",
   42184 => x"208208",
   42185 => x"208208",
   42186 => x"208208",
   42187 => x"208208",
   42188 => x"208208",
   42189 => x"208208",
   42190 => x"208208",
   42191 => x"208208",
   42192 => x"208208",
   42193 => x"208208",
   42194 => x"208208",
   42195 => x"208104",
   42196 => x"104104",
   42197 => x"104104",
   42198 => x"104104",
   42199 => x"104104",
   42200 => x"104104",
   42201 => x"104104",
   42202 => x"104104",
   42203 => x"104104",
   42204 => x"104104",
   42205 => x"104104",
   42206 => x"104104",
   42207 => x"104104",
   42208 => x"104104",
   42209 => x"104104",
   42210 => x"104104",
   42211 => x"104104",
   42212 => x"104104",
   42213 => x"104104",
   42214 => x"104104",
   42215 => x"104104",
   42216 => x"104104",
   42217 => x"104104",
   42218 => x"104000",
   42219 => x"000000",
   42220 => x"000000",
   42221 => x"000000",
   42222 => x"000000",
   42223 => x"000000",
   42224 => x"000000",
   42225 => x"000000",
   42226 => x"000000",
   42227 => x"000000",
   42228 => x"000000",
   42229 => x"00057f",
   42230 => x"ffffff",
   42231 => x"ffffff",
   42232 => x"ffffff",
   42233 => x"ffffff",
   42234 => x"ffffff",
   42235 => x"ffffff",
   42236 => x"ffffff",
   42237 => x"ffffff",
   42238 => x"ffffff",
   42239 => x"ffffff",
   42240 => x"ffffff",
   42241 => x"ffffff",
   42242 => x"ffffff",
   42243 => x"ffffff",
   42244 => x"ffffff",
   42245 => x"ffffff",
   42246 => x"ffffff",
   42247 => x"ffffff",
   42248 => x"ffffff",
   42249 => x"ffffff",
   42250 => x"ffffff",
   42251 => x"ffffff",
   42252 => x"ffffff",
   42253 => x"ffffff",
   42254 => x"ffffff",
   42255 => x"ffffff",
   42256 => x"ffffff",
   42257 => x"ffffff",
   42258 => x"ffffff",
   42259 => x"ffffff",
   42260 => x"5c30c3",
   42261 => x"0c30c3",
   42262 => x"0c30c3",
   42263 => x"0c30c3",
   42264 => x"0c30c3",
   42265 => x"0c30c3",
   42266 => x"0c30c3",
   42267 => x"0c30c3",
   42268 => x"0c30c3",
   42269 => x"0c30c3",
   42270 => x"0c30c3",
   42271 => x"0c30c3",
   42272 => x"0c30c3",
   42273 => x"0c30c3",
   42274 => x"0c30c3",
   42275 => x"0c30c3",
   42276 => x"0c30c3",
   42277 => x"0c30c3",
   42278 => x"0c30c3",
   42279 => x"0c30c3",
   42280 => x"0c30c3",
   42281 => x"0c30c3",
   42282 => x"0c30c3",
   42283 => x"0c30c3",
   42284 => x"0c30c3",
   42285 => x"0c30c3",
   42286 => x"0c30c3",
   42287 => x"0c30c3",
   42288 => x"0c3aff",
   42289 => x"ffffff",
   42290 => x"ffffff",
   42291 => x"fffa80",
   42292 => x"00003f",
   42293 => x"ffffff",
   42294 => x"ffffff",
   42295 => x"fff540",
   42296 => x"00057f",
   42297 => x"ffffff",
   42298 => x"ffffff",
   42299 => x"ffffff",
   42300 => x"ffffff",
   42301 => x"ffffff",
   42302 => x"ffffff",
   42303 => x"ffffff",
   42304 => x"ffffff",
   42305 => x"ffffff",
   42306 => x"ffffff",
   42307 => x"ffffff",
   42308 => x"ffffff",
   42309 => x"fffa95",
   42310 => x"abffff",
   42311 => x"ffffff",
   42312 => x"ffffff",
   42313 => x"ffffff",
   42314 => x"ffffff",
   42315 => x"ffffff",
   42316 => x"ffffff",
   42317 => x"ffffff",
   42318 => x"ffffff",
   42319 => x"ffffff",
   42320 => x"ffffff",
   42321 => x"fffb8c",
   42322 => x"30c30c",
   42323 => x"30c30c",
   42324 => x"30c30c",
   42325 => x"30c30c",
   42326 => x"30c30c",
   42327 => x"30c30c",
   42328 => x"30c30c",
   42329 => x"30c30c",
   42330 => x"30c30c",
   42331 => x"30c30c",
   42332 => x"30c30c",
   42333 => x"208208",
   42334 => x"208208",
   42335 => x"208208",
   42336 => x"208208",
   42337 => x"208208",
   42338 => x"208208",
   42339 => x"208208",
   42340 => x"208208",
   42341 => x"208208",
   42342 => x"208208",
   42343 => x"208208",
   42344 => x"208208",
   42345 => x"208208",
   42346 => x"208208",
   42347 => x"208208",
   42348 => x"208208",
   42349 => x"208208",
   42350 => x"208208",
   42351 => x"208208",
   42352 => x"208208",
   42353 => x"208208",
   42354 => x"208208",
   42355 => x"208104",
   42356 => x"104104",
   42357 => x"104104",
   42358 => x"104104",
   42359 => x"104104",
   42360 => x"104104",
   42361 => x"104104",
   42362 => x"104104",
   42363 => x"104104",
   42364 => x"104104",
   42365 => x"104104",
   42366 => x"104104",
   42367 => x"104104",
   42368 => x"104104",
   42369 => x"104104",
   42370 => x"104104",
   42371 => x"104104",
   42372 => x"104104",
   42373 => x"104104",
   42374 => x"104104",
   42375 => x"104104",
   42376 => x"104104",
   42377 => x"104104",
   42378 => x"104000",
   42379 => x"000000",
   42380 => x"000000",
   42381 => x"000000",
   42382 => x"000000",
   42383 => x"000000",
   42384 => x"000000",
   42385 => x"000000",
   42386 => x"000000",
   42387 => x"000000",
   42388 => x"000000",
   42389 => x"00057f",
   42390 => x"ffffff",
   42391 => x"ffffff",
   42392 => x"ffffff",
   42393 => x"ffffff",
   42394 => x"ffffff",
   42395 => x"ffffff",
   42396 => x"ffffff",
   42397 => x"ffffff",
   42398 => x"ffffff",
   42399 => x"ffffff",
   42400 => x"ffffff",
   42401 => x"ffffff",
   42402 => x"ffffff",
   42403 => x"ffffff",
   42404 => x"ffffff",
   42405 => x"ffffff",
   42406 => x"ffffff",
   42407 => x"ffffff",
   42408 => x"ffffff",
   42409 => x"ffffff",
   42410 => x"ffffff",
   42411 => x"ffffff",
   42412 => x"ffffff",
   42413 => x"ffffff",
   42414 => x"ffffff",
   42415 => x"ffffff",
   42416 => x"ffffff",
   42417 => x"ffffff",
   42418 => x"ffffff",
   42419 => x"ffffff",
   42420 => x"feb0c3",
   42421 => x"0c30c3",
   42422 => x"0c30c3",
   42423 => x"0c30c3",
   42424 => x"0c30c3",
   42425 => x"0c30c3",
   42426 => x"0c30c3",
   42427 => x"0c30c3",
   42428 => x"0c30c3",
   42429 => x"0c30c3",
   42430 => x"0c30c3",
   42431 => x"0c30c3",
   42432 => x"0c30c3",
   42433 => x"0c30c3",
   42434 => x"0c30c3",
   42435 => x"0c30c3",
   42436 => x"0c30c3",
   42437 => x"0c30c3",
   42438 => x"0c30c3",
   42439 => x"0c30c3",
   42440 => x"0c30c3",
   42441 => x"0c30c3",
   42442 => x"0c30c3",
   42443 => x"0c30c3",
   42444 => x"0c30c3",
   42445 => x"0c30c3",
   42446 => x"0c30c3",
   42447 => x"0c30c3",
   42448 => x"5ebfff",
   42449 => x"ffffff",
   42450 => x"ffffff",
   42451 => x"fffa80",
   42452 => x"00002a",
   42453 => x"ffffff",
   42454 => x"ffffff",
   42455 => x"a95000",
   42456 => x"015abf",
   42457 => x"ffffff",
   42458 => x"ffffff",
   42459 => x"ffffff",
   42460 => x"ffffff",
   42461 => x"ffffff",
   42462 => x"ffffff",
   42463 => x"ffffff",
   42464 => x"ffffff",
   42465 => x"ffffff",
   42466 => x"ffffff",
   42467 => x"ffffff",
   42468 => x"ffffff",
   42469 => x"fffa95",
   42470 => x"abffff",
   42471 => x"ffffff",
   42472 => x"ffffff",
   42473 => x"ffffff",
   42474 => x"ffffff",
   42475 => x"ffffff",
   42476 => x"ffffff",
   42477 => x"ffffff",
   42478 => x"ffffff",
   42479 => x"ffffff",
   42480 => x"ffffff",
   42481 => x"fffb8c",
   42482 => x"30c30c",
   42483 => x"30c30c",
   42484 => x"30c30c",
   42485 => x"30c30c",
   42486 => x"30c30c",
   42487 => x"30c30c",
   42488 => x"30c30c",
   42489 => x"30c30c",
   42490 => x"30c30c",
   42491 => x"30c30c",
   42492 => x"30c30c",
   42493 => x"208208",
   42494 => x"208208",
   42495 => x"208208",
   42496 => x"208208",
   42497 => x"208208",
   42498 => x"208208",
   42499 => x"208208",
   42500 => x"208208",
   42501 => x"208208",
   42502 => x"208208",
   42503 => x"208208",
   42504 => x"208208",
   42505 => x"208208",
   42506 => x"208208",
   42507 => x"208208",
   42508 => x"208208",
   42509 => x"208208",
   42510 => x"208208",
   42511 => x"208208",
   42512 => x"208208",
   42513 => x"208208",
   42514 => x"208208",
   42515 => x"208104",
   42516 => x"104104",
   42517 => x"104104",
   42518 => x"104104",
   42519 => x"104104",
   42520 => x"104104",
   42521 => x"104104",
   42522 => x"104104",
   42523 => x"104104",
   42524 => x"104104",
   42525 => x"104104",
   42526 => x"104104",
   42527 => x"104104",
   42528 => x"104104",
   42529 => x"104104",
   42530 => x"104104",
   42531 => x"104104",
   42532 => x"104104",
   42533 => x"104104",
   42534 => x"104104",
   42535 => x"104104",
   42536 => x"104104",
   42537 => x"104104",
   42538 => x"104000",
   42539 => x"000000",
   42540 => x"000000",
   42541 => x"000000",
   42542 => x"000000",
   42543 => x"000000",
   42544 => x"000000",
   42545 => x"000000",
   42546 => x"000000",
   42547 => x"000000",
   42548 => x"000000",
   42549 => x"00057f",
   42550 => x"ffffff",
   42551 => x"ffffff",
   42552 => x"ffffff",
   42553 => x"ffffff",
   42554 => x"ffffff",
   42555 => x"ffffff",
   42556 => x"ffffff",
   42557 => x"ffffff",
   42558 => x"ffffff",
   42559 => x"ffffff",
   42560 => x"ffffff",
   42561 => x"ffffff",
   42562 => x"ffffff",
   42563 => x"ffffff",
   42564 => x"ffffff",
   42565 => x"ffffff",
   42566 => x"ffffff",
   42567 => x"ffffff",
   42568 => x"ffffff",
   42569 => x"ffffff",
   42570 => x"ffffff",
   42571 => x"ffffff",
   42572 => x"ffffff",
   42573 => x"ffffff",
   42574 => x"ffffff",
   42575 => x"ffffff",
   42576 => x"ffffff",
   42577 => x"ffffff",
   42578 => x"ffffff",
   42579 => x"ffffff",
   42580 => x"fffad7",
   42581 => x"0c30c3",
   42582 => x"0c30c3",
   42583 => x"0c30c3",
   42584 => x"0c30c3",
   42585 => x"0c30c3",
   42586 => x"0c30c3",
   42587 => x"0c30c3",
   42588 => x"0c30c3",
   42589 => x"0c30c3",
   42590 => x"0c30c3",
   42591 => x"0c30c3",
   42592 => x"0c30c3",
   42593 => x"0c30c3",
   42594 => x"0c30c3",
   42595 => x"0c30c3",
   42596 => x"0c30c3",
   42597 => x"0c30c3",
   42598 => x"0c30c3",
   42599 => x"0c30c3",
   42600 => x"0c30c3",
   42601 => x"0c30c3",
   42602 => x"0c30c3",
   42603 => x"0c30c3",
   42604 => x"0c30c3",
   42605 => x"0c30c3",
   42606 => x"0c30c3",
   42607 => x"0c30d7",
   42608 => x"afffff",
   42609 => x"ffffff",
   42610 => x"ffffff",
   42611 => x"fffa80",
   42612 => x"000015",
   42613 => x"555555",
   42614 => x"555555",
   42615 => x"000000",
   42616 => x"56afff",
   42617 => x"ffffff",
   42618 => x"ffffff",
   42619 => x"ffffff",
   42620 => x"ffffff",
   42621 => x"ffffff",
   42622 => x"ffffff",
   42623 => x"ffffff",
   42624 => x"ffffff",
   42625 => x"ffffff",
   42626 => x"ffffff",
   42627 => x"ffffff",
   42628 => x"ffffff",
   42629 => x"fffa95",
   42630 => x"abffff",
   42631 => x"ffffff",
   42632 => x"ffffff",
   42633 => x"ffffff",
   42634 => x"ffffff",
   42635 => x"ffffff",
   42636 => x"ffffff",
   42637 => x"ffffff",
   42638 => x"ffffff",
   42639 => x"ffffff",
   42640 => x"ffffff",
   42641 => x"fffb8c",
   42642 => x"30c30c",
   42643 => x"30c30c",
   42644 => x"30c30c",
   42645 => x"30c30c",
   42646 => x"30c30c",
   42647 => x"30c30c",
   42648 => x"30c30c",
   42649 => x"30c30c",
   42650 => x"30c30c",
   42651 => x"30c30c",
   42652 => x"30c30c",
   42653 => x"208208",
   42654 => x"208208",
   42655 => x"208208",
   42656 => x"208208",
   42657 => x"208208",
   42658 => x"208208",
   42659 => x"208208",
   42660 => x"208208",
   42661 => x"208208",
   42662 => x"208208",
   42663 => x"208208",
   42664 => x"208208",
   42665 => x"208208",
   42666 => x"208208",
   42667 => x"208208",
   42668 => x"208208",
   42669 => x"208208",
   42670 => x"208208",
   42671 => x"208208",
   42672 => x"208208",
   42673 => x"208208",
   42674 => x"208208",
   42675 => x"208104",
   42676 => x"104104",
   42677 => x"104104",
   42678 => x"104104",
   42679 => x"104104",
   42680 => x"104104",
   42681 => x"104104",
   42682 => x"104104",
   42683 => x"104104",
   42684 => x"104104",
   42685 => x"104104",
   42686 => x"104104",
   42687 => x"104104",
   42688 => x"104104",
   42689 => x"104104",
   42690 => x"104104",
   42691 => x"104104",
   42692 => x"104104",
   42693 => x"104104",
   42694 => x"104104",
   42695 => x"104104",
   42696 => x"104104",
   42697 => x"104104",
   42698 => x"104000",
   42699 => x"000000",
   42700 => x"000000",
   42701 => x"000000",
   42702 => x"000000",
   42703 => x"000000",
   42704 => x"000000",
   42705 => x"000000",
   42706 => x"000000",
   42707 => x"000000",
   42708 => x"000000",
   42709 => x"00057f",
   42710 => x"ffffff",
   42711 => x"ffffff",
   42712 => x"ffffff",
   42713 => x"ffffff",
   42714 => x"ffffff",
   42715 => x"ffffff",
   42716 => x"ffffff",
   42717 => x"ffffff",
   42718 => x"ffffff",
   42719 => x"ffffff",
   42720 => x"ffffff",
   42721 => x"ffffff",
   42722 => x"ffffff",
   42723 => x"ffffff",
   42724 => x"ffffff",
   42725 => x"ffffff",
   42726 => x"ffffff",
   42727 => x"ffffff",
   42728 => x"ffffff",
   42729 => x"ffffff",
   42730 => x"ffffff",
   42731 => x"ffffff",
   42732 => x"ffffff",
   42733 => x"ffffff",
   42734 => x"ffffff",
   42735 => x"ffffff",
   42736 => x"ffffff",
   42737 => x"ffffff",
   42738 => x"ffffff",
   42739 => x"ffffff",
   42740 => x"ffffeb",
   42741 => x"5c30c3",
   42742 => x"0c30c3",
   42743 => x"0c30c3",
   42744 => x"0c30c3",
   42745 => x"0c30c3",
   42746 => x"0c30c3",
   42747 => x"0c30c3",
   42748 => x"0c30c3",
   42749 => x"0c30c3",
   42750 => x"0c30c3",
   42751 => x"0c30c3",
   42752 => x"0c30c3",
   42753 => x"0c30c3",
   42754 => x"0c30c3",
   42755 => x"0c30c3",
   42756 => x"0c30c3",
   42757 => x"0c30c3",
   42758 => x"0c30c3",
   42759 => x"0c30c3",
   42760 => x"0c30c3",
   42761 => x"0c30c3",
   42762 => x"0c30c3",
   42763 => x"0c30c3",
   42764 => x"0c30c3",
   42765 => x"0c30c3",
   42766 => x"0c30c3",
   42767 => x"0c3aff",
   42768 => x"ffffff",
   42769 => x"ffffff",
   42770 => x"ffffff",
   42771 => x"fffa80",
   42772 => x"000000",
   42773 => x"000000",
   42774 => x"000000",
   42775 => x"00056a",
   42776 => x"abffff",
   42777 => x"ffffff",
   42778 => x"ffffff",
   42779 => x"ffffff",
   42780 => x"ffffff",
   42781 => x"ffffff",
   42782 => x"ffffff",
   42783 => x"ffffff",
   42784 => x"ffffff",
   42785 => x"ffffff",
   42786 => x"ffffff",
   42787 => x"ffffff",
   42788 => x"ffffff",
   42789 => x"fffa95",
   42790 => x"abffff",
   42791 => x"ffffff",
   42792 => x"ffffff",
   42793 => x"ffffff",
   42794 => x"ffffff",
   42795 => x"ffffff",
   42796 => x"ffffff",
   42797 => x"ffffff",
   42798 => x"ffffff",
   42799 => x"ffffff",
   42800 => x"ffffff",
   42801 => x"fffb8c",
   42802 => x"30c30c",
   42803 => x"30c30c",
   42804 => x"30c30c",
   42805 => x"30c30c",
   42806 => x"30c30c",
   42807 => x"30c30c",
   42808 => x"30c30c",
   42809 => x"30c30c",
   42810 => x"30c30c",
   42811 => x"30c30c",
   42812 => x"30c30c",
   42813 => x"208208",
   42814 => x"208208",
   42815 => x"208208",
   42816 => x"208208",
   42817 => x"208208",
   42818 => x"208208",
   42819 => x"208208",
   42820 => x"208208",
   42821 => x"208208",
   42822 => x"208208",
   42823 => x"208208",
   42824 => x"208208",
   42825 => x"208208",
   42826 => x"208208",
   42827 => x"208208",
   42828 => x"208208",
   42829 => x"208208",
   42830 => x"208208",
   42831 => x"208208",
   42832 => x"208208",
   42833 => x"208208",
   42834 => x"208208",
   42835 => x"208104",
   42836 => x"104104",
   42837 => x"104104",
   42838 => x"104104",
   42839 => x"104104",
   42840 => x"104104",
   42841 => x"104104",
   42842 => x"104104",
   42843 => x"104104",
   42844 => x"104104",
   42845 => x"104104",
   42846 => x"104104",
   42847 => x"104104",
   42848 => x"104104",
   42849 => x"104104",
   42850 => x"104104",
   42851 => x"104104",
   42852 => x"104104",
   42853 => x"104104",
   42854 => x"104104",
   42855 => x"104104",
   42856 => x"104104",
   42857 => x"104104",
   42858 => x"104000",
   42859 => x"000000",
   42860 => x"000000",
   42861 => x"000000",
   42862 => x"000000",
   42863 => x"000000",
   42864 => x"000000",
   42865 => x"000000",
   42866 => x"000000",
   42867 => x"000000",
   42868 => x"000000",
   42869 => x"00057f",
   42870 => x"ffffff",
   42871 => x"ffffff",
   42872 => x"ffffff",
   42873 => x"ffffff",
   42874 => x"ffffff",
   42875 => x"ffffff",
   42876 => x"ffffff",
   42877 => x"ffffff",
   42878 => x"ffffff",
   42879 => x"ffffff",
   42880 => x"ffffff",
   42881 => x"ffffff",
   42882 => x"ffffff",
   42883 => x"ffffff",
   42884 => x"ffffff",
   42885 => x"ffffff",
   42886 => x"ffffff",
   42887 => x"ffffff",
   42888 => x"ffffff",
   42889 => x"ffffff",
   42890 => x"ffffff",
   42891 => x"ffffff",
   42892 => x"ffffff",
   42893 => x"ffffff",
   42894 => x"ffffff",
   42895 => x"ffffff",
   42896 => x"ffffff",
   42897 => x"ffffff",
   42898 => x"ffffff",
   42899 => x"ffffff",
   42900 => x"ffffff",
   42901 => x"feb0c3",
   42902 => x"0c30c3",
   42903 => x"0c30c3",
   42904 => x"0c30c3",
   42905 => x"0c30c3",
   42906 => x"0c30c3",
   42907 => x"0c30c3",
   42908 => x"0c30c3",
   42909 => x"0c30c3",
   42910 => x"0c30c3",
   42911 => x"0c30c3",
   42912 => x"0c30c3",
   42913 => x"0c30c3",
   42914 => x"0c30c3",
   42915 => x"0c30c3",
   42916 => x"0c30c3",
   42917 => x"0c30c3",
   42918 => x"0c30c3",
   42919 => x"0c30c3",
   42920 => x"0c30c3",
   42921 => x"0c30c3",
   42922 => x"0c30c3",
   42923 => x"0c30c3",
   42924 => x"0c30c3",
   42925 => x"0c30c3",
   42926 => x"0c30c3",
   42927 => x"5ebfff",
   42928 => x"ffffff",
   42929 => x"ffffff",
   42930 => x"ffffff",
   42931 => x"fffa80",
   42932 => x"000000",
   42933 => x"000000",
   42934 => x"000000",
   42935 => x"000015",
   42936 => x"abffff",
   42937 => x"ffffff",
   42938 => x"ffffff",
   42939 => x"ffffff",
   42940 => x"ffffff",
   42941 => x"ffffff",
   42942 => x"ffffff",
   42943 => x"ffffff",
   42944 => x"ffffff",
   42945 => x"ffffff",
   42946 => x"ffffff",
   42947 => x"ffffff",
   42948 => x"ffffff",
   42949 => x"fffa95",
   42950 => x"abffff",
   42951 => x"ffffff",
   42952 => x"ffffff",
   42953 => x"ffffff",
   42954 => x"ffffff",
   42955 => x"ffffff",
   42956 => x"ffffff",
   42957 => x"ffffff",
   42958 => x"ffffff",
   42959 => x"ffffff",
   42960 => x"ffffff",
   42961 => x"fffb8c",
   42962 => x"30c30c",
   42963 => x"30c30c",
   42964 => x"30c30c",
   42965 => x"30c30c",
   42966 => x"30c30c",
   42967 => x"30c30c",
   42968 => x"30c30c",
   42969 => x"30c30c",
   42970 => x"30c30c",
   42971 => x"30c30c",
   42972 => x"30c30c",
   42973 => x"208208",
   42974 => x"208208",
   42975 => x"208208",
   42976 => x"208208",
   42977 => x"208208",
   42978 => x"208208",
   42979 => x"208208",
   42980 => x"208208",
   42981 => x"208208",
   42982 => x"208208",
   42983 => x"208208",
   42984 => x"208208",
   42985 => x"208208",
   42986 => x"208208",
   42987 => x"208208",
   42988 => x"208208",
   42989 => x"208208",
   42990 => x"208208",
   42991 => x"208208",
   42992 => x"208208",
   42993 => x"208208",
   42994 => x"208208",
   42995 => x"208104",
   42996 => x"104104",
   42997 => x"104104",
   42998 => x"104104",
   42999 => x"104104",
   43000 => x"104104",
   43001 => x"104104",
   43002 => x"104104",
   43003 => x"104104",
   43004 => x"104104",
   43005 => x"104104",
   43006 => x"104104",
   43007 => x"104104",
   43008 => x"104104",
   43009 => x"104104",
   43010 => x"104104",
   43011 => x"104104",
   43012 => x"104104",
   43013 => x"104104",
   43014 => x"104104",
   43015 => x"104104",
   43016 => x"104104",
   43017 => x"104104",
   43018 => x"104000",
   43019 => x"000000",
   43020 => x"000000",
   43021 => x"000000",
   43022 => x"000000",
   43023 => x"000000",
   43024 => x"000000",
   43025 => x"000000",
   43026 => x"000000",
   43027 => x"000000",
   43028 => x"000000",
   43029 => x"00057f",
   43030 => x"ffffff",
   43031 => x"ffffff",
   43032 => x"ffffff",
   43033 => x"ffffff",
   43034 => x"ffffff",
   43035 => x"ffffff",
   43036 => x"ffffff",
   43037 => x"ffffff",
   43038 => x"ffffff",
   43039 => x"ffffff",
   43040 => x"ffffff",
   43041 => x"ffffff",
   43042 => x"ffffff",
   43043 => x"ffffff",
   43044 => x"ffffff",
   43045 => x"ffffff",
   43046 => x"ffffff",
   43047 => x"ffffff",
   43048 => x"ffffff",
   43049 => x"ffffff",
   43050 => x"ffffff",
   43051 => x"ffffff",
   43052 => x"ffffff",
   43053 => x"ffffff",
   43054 => x"ffffff",
   43055 => x"ffffff",
   43056 => x"ffffff",
   43057 => x"ffffff",
   43058 => x"ffffff",
   43059 => x"ffffff",
   43060 => x"ffffff",
   43061 => x"fffad7",
   43062 => x"0c30c3",
   43063 => x"0c30c3",
   43064 => x"0c30c3",
   43065 => x"0c30c3",
   43066 => x"0c30c3",
   43067 => x"0c30c3",
   43068 => x"0c30c3",
   43069 => x"0c30c3",
   43070 => x"0c30c3",
   43071 => x"0c30c3",
   43072 => x"0c30c3",
   43073 => x"0c30c3",
   43074 => x"0c30c3",
   43075 => x"0c30c3",
   43076 => x"0c30c3",
   43077 => x"0c30c3",
   43078 => x"0c30c3",
   43079 => x"0c30c3",
   43080 => x"0c30c3",
   43081 => x"0c30c3",
   43082 => x"0c30c3",
   43083 => x"0c30c3",
   43084 => x"0c30c3",
   43085 => x"0c30c3",
   43086 => x"0c30eb",
   43087 => x"ffffff",
   43088 => x"ffffff",
   43089 => x"ffffff",
   43090 => x"ffffff",
   43091 => x"fffa80",
   43092 => x"000015",
   43093 => x"555555",
   43094 => x"555540",
   43095 => x"000000",
   43096 => x"56afff",
   43097 => x"ffffff",
   43098 => x"ffffff",
   43099 => x"ffffff",
   43100 => x"ffffff",
   43101 => x"ffffff",
   43102 => x"ffffff",
   43103 => x"ffffff",
   43104 => x"ffffff",
   43105 => x"ffffff",
   43106 => x"ffffff",
   43107 => x"ffffff",
   43108 => x"ffffff",
   43109 => x"fffa95",
   43110 => x"abffff",
   43111 => x"ffffff",
   43112 => x"ffffff",
   43113 => x"ffffff",
   43114 => x"ffffff",
   43115 => x"ffffff",
   43116 => x"ffffff",
   43117 => x"ffffff",
   43118 => x"ffffff",
   43119 => x"ffffff",
   43120 => x"ffffff",
   43121 => x"fffb8c",
   43122 => x"30c30c",
   43123 => x"30c30c",
   43124 => x"30c30c",
   43125 => x"30c30c",
   43126 => x"30c30c",
   43127 => x"30c30c",
   43128 => x"30c30c",
   43129 => x"30c30c",
   43130 => x"30c30c",
   43131 => x"30c30c",
   43132 => x"30c30c",
   43133 => x"208208",
   43134 => x"208208",
   43135 => x"208208",
   43136 => x"208208",
   43137 => x"208208",
   43138 => x"208208",
   43139 => x"208208",
   43140 => x"208208",
   43141 => x"208208",
   43142 => x"208208",
   43143 => x"208208",
   43144 => x"208208",
   43145 => x"208208",
   43146 => x"208208",
   43147 => x"208208",
   43148 => x"208208",
   43149 => x"208208",
   43150 => x"208208",
   43151 => x"208208",
   43152 => x"208208",
   43153 => x"208208",
   43154 => x"208208",
   43155 => x"208104",
   43156 => x"104104",
   43157 => x"104104",
   43158 => x"104104",
   43159 => x"104104",
   43160 => x"104104",
   43161 => x"104104",
   43162 => x"104104",
   43163 => x"104104",
   43164 => x"104104",
   43165 => x"104104",
   43166 => x"104104",
   43167 => x"104104",
   43168 => x"104104",
   43169 => x"104104",
   43170 => x"104104",
   43171 => x"104104",
   43172 => x"104104",
   43173 => x"104104",
   43174 => x"104104",
   43175 => x"104104",
   43176 => x"104104",
   43177 => x"104104",
   43178 => x"104000",
   43179 => x"000000",
   43180 => x"000000",
   43181 => x"000000",
   43182 => x"000000",
   43183 => x"000000",
   43184 => x"000000",
   43185 => x"000000",
   43186 => x"000000",
   43187 => x"000000",
   43188 => x"000000",
   43189 => x"00057f",
   43190 => x"ffffff",
   43191 => x"ffffff",
   43192 => x"ffffff",
   43193 => x"ffffff",
   43194 => x"ffffff",
   43195 => x"ffffff",
   43196 => x"ffffff",
   43197 => x"ffffff",
   43198 => x"ffffff",
   43199 => x"ffffff",
   43200 => x"ffffff",
   43201 => x"ffffff",
   43202 => x"ffffff",
   43203 => x"ffffff",
   43204 => x"ffffff",
   43205 => x"ffffff",
   43206 => x"ffffff",
   43207 => x"ffffff",
   43208 => x"ffffff",
   43209 => x"ffffff",
   43210 => x"ffffff",
   43211 => x"ffffff",
   43212 => x"ffffff",
   43213 => x"ffffff",
   43214 => x"ffffff",
   43215 => x"ffffff",
   43216 => x"ffffff",
   43217 => x"ffffff",
   43218 => x"ffffff",
   43219 => x"ffffff",
   43220 => x"ffffff",
   43221 => x"ffffff",
   43222 => x"ad70c3",
   43223 => x"0c30c3",
   43224 => x"0c30c3",
   43225 => x"0c30c3",
   43226 => x"0c30c3",
   43227 => x"0c30c3",
   43228 => x"0c30c3",
   43229 => x"0c30c3",
   43230 => x"0c30c3",
   43231 => x"0c30c3",
   43232 => x"0c30c3",
   43233 => x"0c30c3",
   43234 => x"0c30c3",
   43235 => x"0c30c3",
   43236 => x"0c30c3",
   43237 => x"0c30c3",
   43238 => x"0c30c3",
   43239 => x"0c30c3",
   43240 => x"0c30c3",
   43241 => x"0c30c3",
   43242 => x"0c30c3",
   43243 => x"0c30c3",
   43244 => x"0c30c3",
   43245 => x"0c30c3",
   43246 => x"0d7aff",
   43247 => x"ffffff",
   43248 => x"ffffff",
   43249 => x"ffffff",
   43250 => x"ffffff",
   43251 => x"fffa80",
   43252 => x"00002a",
   43253 => x"ffffff",
   43254 => x"fffaaa",
   43255 => x"a95000",
   43256 => x"00057f",
   43257 => x"ffffff",
   43258 => x"ffffff",
   43259 => x"ffffff",
   43260 => x"ffffff",
   43261 => x"ffffff",
   43262 => x"ffffff",
   43263 => x"ffffff",
   43264 => x"ffffff",
   43265 => x"ffffff",
   43266 => x"ffffff",
   43267 => x"ffffff",
   43268 => x"ffffff",
   43269 => x"fffa95",
   43270 => x"abffff",
   43271 => x"ffffff",
   43272 => x"ffffff",
   43273 => x"ffffff",
   43274 => x"ffffff",
   43275 => x"ffffff",
   43276 => x"ffffff",
   43277 => x"ffffff",
   43278 => x"ffffff",
   43279 => x"ffffff",
   43280 => x"ffffff",
   43281 => x"fffb8c",
   43282 => x"30c30c",
   43283 => x"30c30c",
   43284 => x"30c30c",
   43285 => x"30c30c",
   43286 => x"30c30c",
   43287 => x"30c30c",
   43288 => x"30c30c",
   43289 => x"30c30c",
   43290 => x"30c30c",
   43291 => x"30c30c",
   43292 => x"30c30c",
   43293 => x"208208",
   43294 => x"208208",
   43295 => x"208208",
   43296 => x"208208",
   43297 => x"208208",
   43298 => x"208208",
   43299 => x"208208",
   43300 => x"208208",
   43301 => x"208208",
   43302 => x"208208",
   43303 => x"208208",
   43304 => x"208208",
   43305 => x"208208",
   43306 => x"208208",
   43307 => x"208208",
   43308 => x"208208",
   43309 => x"208208",
   43310 => x"208208",
   43311 => x"208208",
   43312 => x"208208",
   43313 => x"208208",
   43314 => x"208208",
   43315 => x"208104",
   43316 => x"104104",
   43317 => x"104104",
   43318 => x"104104",
   43319 => x"104104",
   43320 => x"104104",
   43321 => x"104104",
   43322 => x"104104",
   43323 => x"104104",
   43324 => x"104104",
   43325 => x"104104",
   43326 => x"104104",
   43327 => x"104104",
   43328 => x"104104",
   43329 => x"104104",
   43330 => x"104104",
   43331 => x"104104",
   43332 => x"104104",
   43333 => x"104104",
   43334 => x"104104",
   43335 => x"104104",
   43336 => x"104104",
   43337 => x"104104",
   43338 => x"104000",
   43339 => x"000000",
   43340 => x"000000",
   43341 => x"000000",
   43342 => x"000000",
   43343 => x"000000",
   43344 => x"000000",
   43345 => x"000000",
   43346 => x"000000",
   43347 => x"000000",
   43348 => x"000000",
   43349 => x"00057f",
   43350 => x"ffffff",
   43351 => x"ffffff",
   43352 => x"ffffff",
   43353 => x"ffffff",
   43354 => x"ffffff",
   43355 => x"ffffff",
   43356 => x"ffffff",
   43357 => x"ffffff",
   43358 => x"ffffff",
   43359 => x"ffffff",
   43360 => x"ffffff",
   43361 => x"ffffff",
   43362 => x"ffffff",
   43363 => x"ffffff",
   43364 => x"ffffff",
   43365 => x"ffffff",
   43366 => x"ffffff",
   43367 => x"ffffff",
   43368 => x"ffffff",
   43369 => x"ffffff",
   43370 => x"ffffff",
   43371 => x"ffffff",
   43372 => x"ffffff",
   43373 => x"ffffff",
   43374 => x"ffffff",
   43375 => x"ffffff",
   43376 => x"ffffff",
   43377 => x"ffffff",
   43378 => x"ffffff",
   43379 => x"ffffff",
   43380 => x"ffffff",
   43381 => x"ffffff",
   43382 => x"febac3",
   43383 => x"0c30c3",
   43384 => x"0c30c3",
   43385 => x"0c30c3",
   43386 => x"0c30c3",
   43387 => x"0c30c3",
   43388 => x"0c30c3",
   43389 => x"0c30c3",
   43390 => x"0c30c3",
   43391 => x"0c30c3",
   43392 => x"0c30c3",
   43393 => x"0c30c3",
   43394 => x"0c30c3",
   43395 => x"0c30c3",
   43396 => x"0c30c3",
   43397 => x"0c30c3",
   43398 => x"0c30c3",
   43399 => x"0c30c3",
   43400 => x"0c30c3",
   43401 => x"0c30c3",
   43402 => x"0c30c3",
   43403 => x"0c30c3",
   43404 => x"0c30c3",
   43405 => x"0c30d7",
   43406 => x"afffff",
   43407 => x"ffffff",
   43408 => x"ffffff",
   43409 => x"ffffff",
   43410 => x"ffffff",
   43411 => x"fffa80",
   43412 => x"00003f",
   43413 => x"ffffff",
   43414 => x"ffffff",
   43415 => x"fffa80",
   43416 => x"00002a",
   43417 => x"ffffff",
   43418 => x"ffffff",
   43419 => x"ffffff",
   43420 => x"ffffff",
   43421 => x"ffffff",
   43422 => x"ffffff",
   43423 => x"ffffff",
   43424 => x"ffffff",
   43425 => x"ffffff",
   43426 => x"ffffff",
   43427 => x"ffffff",
   43428 => x"ffffff",
   43429 => x"fffa95",
   43430 => x"abffff",
   43431 => x"ffffff",
   43432 => x"ffffff",
   43433 => x"ffffff",
   43434 => x"ffffff",
   43435 => x"ffffff",
   43436 => x"ffffff",
   43437 => x"ffffff",
   43438 => x"ffffff",
   43439 => x"ffffff",
   43440 => x"ffffff",
   43441 => x"fffb8c",
   43442 => x"30c30c",
   43443 => x"30c30c",
   43444 => x"30c30c",
   43445 => x"30c30c",
   43446 => x"30c30c",
   43447 => x"30c30c",
   43448 => x"30c30c",
   43449 => x"30c30c",
   43450 => x"30c30c",
   43451 => x"30c30c",
   43452 => x"30c30c",
   43453 => x"208208",
   43454 => x"208208",
   43455 => x"208208",
   43456 => x"208208",
   43457 => x"208208",
   43458 => x"208208",
   43459 => x"208208",
   43460 => x"208208",
   43461 => x"208208",
   43462 => x"208208",
   43463 => x"208208",
   43464 => x"208208",
   43465 => x"208208",
   43466 => x"208208",
   43467 => x"208208",
   43468 => x"208208",
   43469 => x"208208",
   43470 => x"208208",
   43471 => x"208208",
   43472 => x"208208",
   43473 => x"208208",
   43474 => x"208208",
   43475 => x"208104",
   43476 => x"104104",
   43477 => x"104104",
   43478 => x"104104",
   43479 => x"104104",
   43480 => x"104104",
   43481 => x"104104",
   43482 => x"104104",
   43483 => x"104104",
   43484 => x"104104",
   43485 => x"104104",
   43486 => x"104104",
   43487 => x"104104",
   43488 => x"104104",
   43489 => x"104104",
   43490 => x"104104",
   43491 => x"104104",
   43492 => x"104104",
   43493 => x"104104",
   43494 => x"104104",
   43495 => x"104104",
   43496 => x"104104",
   43497 => x"104104",
   43498 => x"104000",
   43499 => x"000000",
   43500 => x"000000",
   43501 => x"000000",
   43502 => x"000000",
   43503 => x"000000",
   43504 => x"000000",
   43505 => x"000000",
   43506 => x"000000",
   43507 => x"000000",
   43508 => x"000000",
   43509 => x"00057f",
   43510 => x"ffffff",
   43511 => x"ffffff",
   43512 => x"ffffff",
   43513 => x"ffffff",
   43514 => x"ffffff",
   43515 => x"ffffff",
   43516 => x"ffffff",
   43517 => x"ffffff",
   43518 => x"ffffff",
   43519 => x"ffffff",
   43520 => x"ffffff",
   43521 => x"ffffff",
   43522 => x"ffffff",
   43523 => x"ffffff",
   43524 => x"ffffff",
   43525 => x"ffffff",
   43526 => x"ffffff",
   43527 => x"ffffff",
   43528 => x"ffffff",
   43529 => x"ffffff",
   43530 => x"ffffff",
   43531 => x"ffffff",
   43532 => x"ffffff",
   43533 => x"ffffff",
   43534 => x"ffffff",
   43535 => x"ffffff",
   43536 => x"ffffff",
   43537 => x"ffffff",
   43538 => x"ffffff",
   43539 => x"ffffff",
   43540 => x"ffffff",
   43541 => x"ffffff",
   43542 => x"ffffeb",
   43543 => x"5c30c3",
   43544 => x"0c30c3",
   43545 => x"0c30c3",
   43546 => x"0c30c3",
   43547 => x"0c30c3",
   43548 => x"0c30c3",
   43549 => x"0c30c3",
   43550 => x"0c30c3",
   43551 => x"0c30c3",
   43552 => x"0c30c3",
   43553 => x"0c30c3",
   43554 => x"0c30c3",
   43555 => x"0c30c3",
   43556 => x"0c30c3",
   43557 => x"0c30c3",
   43558 => x"0c30c3",
   43559 => x"0c30c3",
   43560 => x"0c30c3",
   43561 => x"0c30c3",
   43562 => x"0c30c3",
   43563 => x"0c30c3",
   43564 => x"0c30c3",
   43565 => x"0c3aeb",
   43566 => x"ffffff",
   43567 => x"ffffff",
   43568 => x"ffffff",
   43569 => x"ffffff",
   43570 => x"ffffff",
   43571 => x"fffa80",
   43572 => x"00003f",
   43573 => x"ffffff",
   43574 => x"ffffff",
   43575 => x"ffffd5",
   43576 => x"000015",
   43577 => x"ffffff",
   43578 => x"ffffff",
   43579 => x"ffffff",
   43580 => x"ffffff",
   43581 => x"ffffff",
   43582 => x"ffffff",
   43583 => x"ffffff",
   43584 => x"ffffff",
   43585 => x"ffffff",
   43586 => x"ffffff",
   43587 => x"ffffff",
   43588 => x"ffffff",
   43589 => x"fffa95",
   43590 => x"abffff",
   43591 => x"ffffff",
   43592 => x"ffffff",
   43593 => x"ffffff",
   43594 => x"ffffff",
   43595 => x"ffffff",
   43596 => x"ffffff",
   43597 => x"ffffff",
   43598 => x"ffffff",
   43599 => x"ffffff",
   43600 => x"ffffff",
   43601 => x"fffb8c",
   43602 => x"30c30c",
   43603 => x"30c30c",
   43604 => x"30c30c",
   43605 => x"30c30c",
   43606 => x"30c30c",
   43607 => x"30c30c",
   43608 => x"30c30c",
   43609 => x"30c30c",
   43610 => x"30c30c",
   43611 => x"30c30c",
   43612 => x"30c30c",
   43613 => x"208208",
   43614 => x"208208",
   43615 => x"208208",
   43616 => x"208208",
   43617 => x"208208",
   43618 => x"208208",
   43619 => x"208208",
   43620 => x"208208",
   43621 => x"208208",
   43622 => x"208208",
   43623 => x"208208",
   43624 => x"208208",
   43625 => x"208208",
   43626 => x"208208",
   43627 => x"208208",
   43628 => x"208208",
   43629 => x"208208",
   43630 => x"208208",
   43631 => x"208208",
   43632 => x"208208",
   43633 => x"208208",
   43634 => x"208208",
   43635 => x"208104",
   43636 => x"104104",
   43637 => x"104104",
   43638 => x"104104",
   43639 => x"104104",
   43640 => x"104104",
   43641 => x"104104",
   43642 => x"104104",
   43643 => x"104104",
   43644 => x"104104",
   43645 => x"104104",
   43646 => x"104104",
   43647 => x"104104",
   43648 => x"104104",
   43649 => x"104104",
   43650 => x"104104",
   43651 => x"104104",
   43652 => x"104104",
   43653 => x"104104",
   43654 => x"104104",
   43655 => x"104104",
   43656 => x"104104",
   43657 => x"104104",
   43658 => x"104000",
   43659 => x"000000",
   43660 => x"000000",
   43661 => x"000000",
   43662 => x"000000",
   43663 => x"000000",
   43664 => x"000000",
   43665 => x"000000",
   43666 => x"000000",
   43667 => x"000000",
   43668 => x"000000",
   43669 => x"00057f",
   43670 => x"ffffff",
   43671 => x"ffffff",
   43672 => x"ffffff",
   43673 => x"ffffff",
   43674 => x"ffffff",
   43675 => x"ffffff",
   43676 => x"ffffff",
   43677 => x"ffffff",
   43678 => x"ffffff",
   43679 => x"ffffff",
   43680 => x"ffffff",
   43681 => x"ffffff",
   43682 => x"ffffff",
   43683 => x"ffffff",
   43684 => x"ffffff",
   43685 => x"ffffff",
   43686 => x"ffffff",
   43687 => x"ffffff",
   43688 => x"ffffff",
   43689 => x"ffffff",
   43690 => x"ffffff",
   43691 => x"ffffff",
   43692 => x"ffffff",
   43693 => x"ffffff",
   43694 => x"ffffff",
   43695 => x"ffffff",
   43696 => x"ffffff",
   43697 => x"ffffff",
   43698 => x"ffffff",
   43699 => x"ffffff",
   43700 => x"ffffff",
   43701 => x"ffffff",
   43702 => x"ffffff",
   43703 => x"feb5c3",
   43704 => x"0c30c3",
   43705 => x"0c30c3",
   43706 => x"0c30c3",
   43707 => x"0c30c3",
   43708 => x"0c30c3",
   43709 => x"0c30c3",
   43710 => x"0c30c3",
   43711 => x"0c30c3",
   43712 => x"0c30c3",
   43713 => x"0c30c3",
   43714 => x"0c30c3",
   43715 => x"0c30c3",
   43716 => x"0c30c3",
   43717 => x"0c30c3",
   43718 => x"0c30c3",
   43719 => x"0c30c3",
   43720 => x"0c30c3",
   43721 => x"0c30c3",
   43722 => x"0c30c3",
   43723 => x"0c30c3",
   43724 => x"0c30d7",
   43725 => x"5ebfff",
   43726 => x"ffffff",
   43727 => x"ffffff",
   43728 => x"ffffff",
   43729 => x"ffffff",
   43730 => x"ffffff",
   43731 => x"fffa80",
   43732 => x"00003f",
   43733 => x"ffffff",
   43734 => x"ffffff",
   43735 => x"ffffea",
   43736 => x"000015",
   43737 => x"abffff",
   43738 => x"ffffff",
   43739 => x"ffffff",
   43740 => x"ffffff",
   43741 => x"ffffff",
   43742 => x"ffffff",
   43743 => x"ffffff",
   43744 => x"ffffff",
   43745 => x"ffffff",
   43746 => x"ffffff",
   43747 => x"ffffff",
   43748 => x"ffffff",
   43749 => x"fffa95",
   43750 => x"abffff",
   43751 => x"ffffff",
   43752 => x"ffffff",
   43753 => x"ffffff",
   43754 => x"ffffff",
   43755 => x"ffffff",
   43756 => x"ffffff",
   43757 => x"ffffff",
   43758 => x"ffffff",
   43759 => x"ffffff",
   43760 => x"ffffff",
   43761 => x"fffb8c",
   43762 => x"30c30c",
   43763 => x"30c30c",
   43764 => x"30c30c",
   43765 => x"30c30c",
   43766 => x"30c30c",
   43767 => x"30c30c",
   43768 => x"30c30c",
   43769 => x"30c30c",
   43770 => x"30c30c",
   43771 => x"30c30c",
   43772 => x"30c30c",
   43773 => x"208208",
   43774 => x"208208",
   43775 => x"208208",
   43776 => x"208208",
   43777 => x"208208",
   43778 => x"208208",
   43779 => x"208208",
   43780 => x"208208",
   43781 => x"208208",
   43782 => x"208208",
   43783 => x"208208",
   43784 => x"208208",
   43785 => x"208208",
   43786 => x"208208",
   43787 => x"208208",
   43788 => x"208208",
   43789 => x"208208",
   43790 => x"208208",
   43791 => x"208208",
   43792 => x"208208",
   43793 => x"208208",
   43794 => x"208208",
   43795 => x"208104",
   43796 => x"104104",
   43797 => x"104104",
   43798 => x"104104",
   43799 => x"104104",
   43800 => x"104104",
   43801 => x"104104",
   43802 => x"104104",
   43803 => x"104104",
   43804 => x"104104",
   43805 => x"104104",
   43806 => x"104104",
   43807 => x"104104",
   43808 => x"104104",
   43809 => x"104104",
   43810 => x"104104",
   43811 => x"104104",
   43812 => x"104104",
   43813 => x"104104",
   43814 => x"104104",
   43815 => x"104104",
   43816 => x"104104",
   43817 => x"104104",
   43818 => x"104000",
   43819 => x"000000",
   43820 => x"000000",
   43821 => x"000000",
   43822 => x"000000",
   43823 => x"000000",
   43824 => x"000000",
   43825 => x"000000",
   43826 => x"000000",
   43827 => x"000000",
   43828 => x"000000",
   43829 => x"00057f",
   43830 => x"ffffff",
   43831 => x"ffffff",
   43832 => x"ffffff",
   43833 => x"ffffff",
   43834 => x"ffffff",
   43835 => x"ffffff",
   43836 => x"ffffff",
   43837 => x"ffffff",
   43838 => x"ffffff",
   43839 => x"ffffff",
   43840 => x"ffffff",
   43841 => x"ffffff",
   43842 => x"ffffff",
   43843 => x"ffffff",
   43844 => x"ffffff",
   43845 => x"ffffff",
   43846 => x"ffffff",
   43847 => x"ffffff",
   43848 => x"ffffff",
   43849 => x"ffffff",
   43850 => x"ffffff",
   43851 => x"ffffff",
   43852 => x"ffffff",
   43853 => x"ffffff",
   43854 => x"ffffff",
   43855 => x"ffffff",
   43856 => x"ffffff",
   43857 => x"ffffff",
   43858 => x"ffffff",
   43859 => x"ffffff",
   43860 => x"ffffff",
   43861 => x"ffffff",
   43862 => x"ffffff",
   43863 => x"ffffeb",
   43864 => x"5c30c3",
   43865 => x"0c30c3",
   43866 => x"0c30c3",
   43867 => x"0c30c3",
   43868 => x"0c30c3",
   43869 => x"0c30c3",
   43870 => x"0c30c3",
   43871 => x"0c30c3",
   43872 => x"0c30c3",
   43873 => x"0c30c3",
   43874 => x"0c30c3",
   43875 => x"0c30c3",
   43876 => x"0c30c3",
   43877 => x"0c30c3",
   43878 => x"0c30c3",
   43879 => x"0c30c3",
   43880 => x"0c30c3",
   43881 => x"0c30c3",
   43882 => x"0c30c3",
   43883 => x"0c30c3",
   43884 => x"0d75eb",
   43885 => x"ffffff",
   43886 => x"ffffff",
   43887 => x"ffffff",
   43888 => x"ffffff",
   43889 => x"ffffff",
   43890 => x"ffffff",
   43891 => x"fffa80",
   43892 => x"00003f",
   43893 => x"ffffff",
   43894 => x"ffffff",
   43895 => x"ffffea",
   43896 => x"540000",
   43897 => x"abffff",
   43898 => x"ffffff",
   43899 => x"ffffff",
   43900 => x"ffffff",
   43901 => x"ffffff",
   43902 => x"ffffff",
   43903 => x"ffffff",
   43904 => x"ffffff",
   43905 => x"ffffff",
   43906 => x"ffffff",
   43907 => x"ffffff",
   43908 => x"ffffff",
   43909 => x"fffa95",
   43910 => x"abffff",
   43911 => x"ffffff",
   43912 => x"ffffff",
   43913 => x"ffffff",
   43914 => x"ffffff",
   43915 => x"ffffff",
   43916 => x"ffffff",
   43917 => x"ffffff",
   43918 => x"ffffff",
   43919 => x"ffffff",
   43920 => x"ffffff",
   43921 => x"fffb8c",
   43922 => x"30c30c",
   43923 => x"30c30c",
   43924 => x"30c30c",
   43925 => x"30c30c",
   43926 => x"30c30c",
   43927 => x"30c30c",
   43928 => x"30c30c",
   43929 => x"30c30c",
   43930 => x"30c30c",
   43931 => x"30c30c",
   43932 => x"30c30c",
   43933 => x"208208",
   43934 => x"208208",
   43935 => x"208208",
   43936 => x"208208",
   43937 => x"208208",
   43938 => x"208208",
   43939 => x"208208",
   43940 => x"208208",
   43941 => x"208208",
   43942 => x"208208",
   43943 => x"208208",
   43944 => x"208208",
   43945 => x"208208",
   43946 => x"208208",
   43947 => x"208208",
   43948 => x"208208",
   43949 => x"208208",
   43950 => x"208208",
   43951 => x"208208",
   43952 => x"208208",
   43953 => x"208208",
   43954 => x"208208",
   43955 => x"208104",
   43956 => x"104104",
   43957 => x"104104",
   43958 => x"104104",
   43959 => x"104104",
   43960 => x"104104",
   43961 => x"104104",
   43962 => x"104104",
   43963 => x"104104",
   43964 => x"104104",
   43965 => x"104104",
   43966 => x"104104",
   43967 => x"104104",
   43968 => x"104104",
   43969 => x"104104",
   43970 => x"104104",
   43971 => x"104104",
   43972 => x"104104",
   43973 => x"104104",
   43974 => x"104104",
   43975 => x"104104",
   43976 => x"104104",
   43977 => x"104104",
   43978 => x"104000",
   43979 => x"000000",
   43980 => x"000000",
   43981 => x"000000",
   43982 => x"000000",
   43983 => x"000000",
   43984 => x"000000",
   43985 => x"000000",
   43986 => x"000000",
   43987 => x"000000",
   43988 => x"000000",
   43989 => x"00057f",
   43990 => x"ffffff",
   43991 => x"ffffff",
   43992 => x"ffffff",
   43993 => x"ffffff",
   43994 => x"ffffff",
   43995 => x"ffffff",
   43996 => x"ffffff",
   43997 => x"ffffff",
   43998 => x"ffffff",
   43999 => x"ffffff",
   44000 => x"ffffff",
   44001 => x"ffffff",
   44002 => x"ffffff",
   44003 => x"ffffff",
   44004 => x"ffffff",
   44005 => x"ffffff",
   44006 => x"ffffff",
   44007 => x"ffffff",
   44008 => x"ffffff",
   44009 => x"ffffff",
   44010 => x"ffffff",
   44011 => x"ffffff",
   44012 => x"ffffff",
   44013 => x"ffffff",
   44014 => x"ffffff",
   44015 => x"ffffff",
   44016 => x"ffffff",
   44017 => x"ffffff",
   44018 => x"ffffff",
   44019 => x"ffffff",
   44020 => x"ffffff",
   44021 => x"ffffff",
   44022 => x"ffffff",
   44023 => x"ffffff",
   44024 => x"feb5c3",
   44025 => x"0c30c3",
   44026 => x"0c30c3",
   44027 => x"0c30c3",
   44028 => x"0c30c3",
   44029 => x"0c30c3",
   44030 => x"0c30c3",
   44031 => x"0c30c3",
   44032 => x"0c30c3",
   44033 => x"0c30c3",
   44034 => x"0c30c3",
   44035 => x"0c30c3",
   44036 => x"0c30c3",
   44037 => x"0c30c3",
   44038 => x"0c30c3",
   44039 => x"0c30c3",
   44040 => x"0c30c3",
   44041 => x"0c30c3",
   44042 => x"0c30c3",
   44043 => x"0c30d7",
   44044 => x"5ebfff",
   44045 => x"ffffff",
   44046 => x"ffffff",
   44047 => x"ffffff",
   44048 => x"ffffff",
   44049 => x"ffffff",
   44050 => x"ffffff",
   44051 => x"fffa80",
   44052 => x"00003f",
   44053 => x"ffffff",
   44054 => x"ffffff",
   44055 => x"ffffea",
   44056 => x"540000",
   44057 => x"abffff",
   44058 => x"ffffff",
   44059 => x"ffffff",
   44060 => x"ffffff",
   44061 => x"ffffff",
   44062 => x"ffffff",
   44063 => x"ffffff",
   44064 => x"ffffff",
   44065 => x"ffffff",
   44066 => x"ffffff",
   44067 => x"ffffff",
   44068 => x"ffffff",
   44069 => x"fffa95",
   44070 => x"abffff",
   44071 => x"ffffff",
   44072 => x"ffffff",
   44073 => x"ffffff",
   44074 => x"ffffff",
   44075 => x"ffffff",
   44076 => x"ffffff",
   44077 => x"ffffff",
   44078 => x"ffffff",
   44079 => x"ffffff",
   44080 => x"ffffff",
   44081 => x"fffb8c",
   44082 => x"30c30c",
   44083 => x"30c30c",
   44084 => x"30c30c",
   44085 => x"30c30c",
   44086 => x"30c30c",
   44087 => x"30c30c",
   44088 => x"30c30c",
   44089 => x"30c30c",
   44090 => x"30c30c",
   44091 => x"30c30c",
   44092 => x"30c30c",
   44093 => x"208208",
   44094 => x"208208",
   44095 => x"208208",
   44096 => x"208208",
   44097 => x"208208",
   44098 => x"208208",
   44099 => x"208208",
   44100 => x"208208",
   44101 => x"208208",
   44102 => x"208208",
   44103 => x"208208",
   44104 => x"208208",
   44105 => x"208208",
   44106 => x"208208",
   44107 => x"208208",
   44108 => x"208208",
   44109 => x"208208",
   44110 => x"208208",
   44111 => x"208208",
   44112 => x"208208",
   44113 => x"208208",
   44114 => x"208208",
   44115 => x"208104",
   44116 => x"104104",
   44117 => x"104104",
   44118 => x"104104",
   44119 => x"104104",
   44120 => x"104104",
   44121 => x"104104",
   44122 => x"104104",
   44123 => x"104104",
   44124 => x"104104",
   44125 => x"104104",
   44126 => x"104104",
   44127 => x"104104",
   44128 => x"104104",
   44129 => x"104104",
   44130 => x"104104",
   44131 => x"104104",
   44132 => x"104104",
   44133 => x"104104",
   44134 => x"104104",
   44135 => x"104104",
   44136 => x"104104",
   44137 => x"104104",
   44138 => x"104000",
   44139 => x"000000",
   44140 => x"000000",
   44141 => x"000000",
   44142 => x"000000",
   44143 => x"000000",
   44144 => x"000000",
   44145 => x"000000",
   44146 => x"000000",
   44147 => x"000000",
   44148 => x"000000",
   44149 => x"00057f",
   44150 => x"ffffff",
   44151 => x"ffffff",
   44152 => x"ffffff",
   44153 => x"ffffff",
   44154 => x"ffffff",
   44155 => x"ffffff",
   44156 => x"ffffff",
   44157 => x"ffffff",
   44158 => x"ffffff",
   44159 => x"ffffff",
   44160 => x"ffffff",
   44161 => x"ffffff",
   44162 => x"ffffff",
   44163 => x"ffffff",
   44164 => x"ffffff",
   44165 => x"ffffff",
   44166 => x"ffffff",
   44167 => x"ffffff",
   44168 => x"ffffff",
   44169 => x"ffffff",
   44170 => x"ffffff",
   44171 => x"ffffff",
   44172 => x"ffffff",
   44173 => x"ffffff",
   44174 => x"ffffff",
   44175 => x"ffffff",
   44176 => x"ffffff",
   44177 => x"ffffff",
   44178 => x"ffffff",
   44179 => x"ffffff",
   44180 => x"ffffff",
   44181 => x"ffffff",
   44182 => x"ffffff",
   44183 => x"ffffff",
   44184 => x"ffffeb",
   44185 => x"5d70c3",
   44186 => x"0c30c3",
   44187 => x"0c30c3",
   44188 => x"0c30c3",
   44189 => x"0c30c3",
   44190 => x"0c30c3",
   44191 => x"0c30c3",
   44192 => x"0c30c3",
   44193 => x"0c30c3",
   44194 => x"0c30c3",
   44195 => x"0c30c3",
   44196 => x"0c30c3",
   44197 => x"0c30c3",
   44198 => x"0c30c3",
   44199 => x"0c30c3",
   44200 => x"0c30c3",
   44201 => x"0c30c3",
   44202 => x"0c30c3",
   44203 => x"0d75eb",
   44204 => x"ffffff",
   44205 => x"ffffff",
   44206 => x"ffffff",
   44207 => x"ffffff",
   44208 => x"ffffff",
   44209 => x"ffffff",
   44210 => x"ffffff",
   44211 => x"fffa80",
   44212 => x"00003f",
   44213 => x"ffffff",
   44214 => x"ffffff",
   44215 => x"ffffea",
   44216 => x"540000",
   44217 => x"abffff",
   44218 => x"ffffff",
   44219 => x"ffffff",
   44220 => x"ffffff",
   44221 => x"ffffff",
   44222 => x"ffffff",
   44223 => x"ffffff",
   44224 => x"ffffff",
   44225 => x"ffffff",
   44226 => x"ffffff",
   44227 => x"ffffff",
   44228 => x"ffffff",
   44229 => x"fffa95",
   44230 => x"abffff",
   44231 => x"ffffff",
   44232 => x"ffffff",
   44233 => x"ffffff",
   44234 => x"ffffff",
   44235 => x"ffffff",
   44236 => x"ffffff",
   44237 => x"ffffff",
   44238 => x"ffffff",
   44239 => x"ffffff",
   44240 => x"ffffff",
   44241 => x"fffb8c",
   44242 => x"30c30c",
   44243 => x"30c30c",
   44244 => x"30c30c",
   44245 => x"30c30c",
   44246 => x"30c30c",
   44247 => x"30c30c",
   44248 => x"30c30c",
   44249 => x"30c30c",
   44250 => x"30c30c",
   44251 => x"30c30c",
   44252 => x"30c30c",
   44253 => x"208208",
   44254 => x"208208",
   44255 => x"208208",
   44256 => x"208208",
   44257 => x"208208",
   44258 => x"208208",
   44259 => x"208208",
   44260 => x"208208",
   44261 => x"208208",
   44262 => x"208208",
   44263 => x"208208",
   44264 => x"208208",
   44265 => x"208208",
   44266 => x"208208",
   44267 => x"208208",
   44268 => x"208208",
   44269 => x"208208",
   44270 => x"208208",
   44271 => x"208208",
   44272 => x"208208",
   44273 => x"208208",
   44274 => x"208208",
   44275 => x"208104",
   44276 => x"104104",
   44277 => x"104104",
   44278 => x"104104",
   44279 => x"104104",
   44280 => x"104104",
   44281 => x"104104",
   44282 => x"104104",
   44283 => x"104104",
   44284 => x"104104",
   44285 => x"104104",
   44286 => x"104104",
   44287 => x"104104",
   44288 => x"104104",
   44289 => x"104104",
   44290 => x"104104",
   44291 => x"104104",
   44292 => x"104104",
   44293 => x"104104",
   44294 => x"104104",
   44295 => x"104104",
   44296 => x"104104",
   44297 => x"104104",
   44298 => x"104000",
   44299 => x"000000",
   44300 => x"000000",
   44301 => x"000000",
   44302 => x"000000",
   44303 => x"000000",
   44304 => x"000000",
   44305 => x"000000",
   44306 => x"000000",
   44307 => x"000000",
   44308 => x"000000",
   44309 => x"00057f",
   44310 => x"ffffff",
   44311 => x"ffffff",
   44312 => x"ffffff",
   44313 => x"ffffff",
   44314 => x"ffffff",
   44315 => x"ffffff",
   44316 => x"ffffff",
   44317 => x"ffffff",
   44318 => x"ffffff",
   44319 => x"ffffff",
   44320 => x"ffffff",
   44321 => x"ffffff",
   44322 => x"ffffff",
   44323 => x"ffffff",
   44324 => x"ffffff",
   44325 => x"ffffff",
   44326 => x"ffffff",
   44327 => x"ffffff",
   44328 => x"ffffff",
   44329 => x"ffffff",
   44330 => x"ffffff",
   44331 => x"ffffff",
   44332 => x"ffffff",
   44333 => x"ffffff",
   44334 => x"ffffff",
   44335 => x"ffffff",
   44336 => x"ffffff",
   44337 => x"ffffff",
   44338 => x"ffffff",
   44339 => x"ffffff",
   44340 => x"ffffff",
   44341 => x"ffffff",
   44342 => x"ffffff",
   44343 => x"ffffff",
   44344 => x"ffffff",
   44345 => x"feb5d7",
   44346 => x"0c30c3",
   44347 => x"0c30c3",
   44348 => x"0c30c3",
   44349 => x"0c30c3",
   44350 => x"0c30c3",
   44351 => x"0c30c3",
   44352 => x"0c30c3",
   44353 => x"0c30c3",
   44354 => x"0c30c3",
   44355 => x"0c30c3",
   44356 => x"0c30c3",
   44357 => x"0c30c3",
   44358 => x"0c30c3",
   44359 => x"0c30c3",
   44360 => x"0c30c3",
   44361 => x"0c30c3",
   44362 => x"0c35d7",
   44363 => x"aebfff",
   44364 => x"ffffff",
   44365 => x"ffffff",
   44366 => x"ffffff",
   44367 => x"ffffff",
   44368 => x"ffffff",
   44369 => x"ffffff",
   44370 => x"ffffff",
   44371 => x"fffa80",
   44372 => x"00003f",
   44373 => x"ffffff",
   44374 => x"ffffff",
   44375 => x"ffffea",
   44376 => x"000000",
   44377 => x"abffff",
   44378 => x"ffffff",
   44379 => x"ffffff",
   44380 => x"ffffff",
   44381 => x"ffffff",
   44382 => x"ffffff",
   44383 => x"ffffff",
   44384 => x"ffffff",
   44385 => x"ffffff",
   44386 => x"ffffff",
   44387 => x"ffffff",
   44388 => x"ffffff",
   44389 => x"fffa95",
   44390 => x"abffff",
   44391 => x"ffffff",
   44392 => x"ffffff",
   44393 => x"ffffff",
   44394 => x"ffffff",
   44395 => x"ffffff",
   44396 => x"ffffff",
   44397 => x"ffffff",
   44398 => x"ffffff",
   44399 => x"ffffff",
   44400 => x"ffffff",
   44401 => x"ffffee",
   44402 => x"75d75d",
   44403 => x"75d75d",
   44404 => x"75d75d",
   44405 => x"75d75d",
   44406 => x"75d75d",
   44407 => x"75d75d",
   44408 => x"75d75d",
   44409 => x"75d75d",
   44410 => x"75d75d",
   44411 => x"75d75d",
   44412 => x"75d75d",
   44413 => x"75d75d",
   44414 => x"75d75d",
   44415 => x"75d75d",
   44416 => x"75d75d",
   44417 => x"75d75d",
   44418 => x"75d75d",
   44419 => x"75d75d",
   44420 => x"75d75d",
   44421 => x"75d75d",
   44422 => x"759659",
   44423 => x"659659",
   44424 => x"659659",
   44425 => x"659659",
   44426 => x"659659",
   44427 => x"659659",
   44428 => x"659659",
   44429 => x"659659",
   44430 => x"659659",
   44431 => x"659659",
   44432 => x"659659",
   44433 => x"659659",
   44434 => x"659659",
   44435 => x"659659",
   44436 => x"659659",
   44437 => x"659659",
   44438 => x"659659",
   44439 => x"659659",
   44440 => x"659659",
   44441 => x"659659",
   44442 => x"659659",
   44443 => x"659659",
   44444 => x"659659",
   44445 => x"659659",
   44446 => x"659659",
   44447 => x"659659",
   44448 => x"659659",
   44449 => x"659659",
   44450 => x"659659",
   44451 => x"659659",
   44452 => x"659659",
   44453 => x"659659",
   44454 => x"659659",
   44455 => x"659659",
   44456 => x"659659",
   44457 => x"659659",
   44458 => x"659659",
   44459 => x"659659",
   44460 => x"659659",
   44461 => x"659659",
   44462 => x"659659",
   44463 => x"659659",
   44464 => x"555555",
   44465 => x"555555",
   44466 => x"555555",
   44467 => x"555555",
   44468 => x"555555",
   44469 => x"555abf",
   44470 => x"ffffff",
   44471 => x"ffffff",
   44472 => x"ffffff",
   44473 => x"ffffff",
   44474 => x"ffffff",
   44475 => x"ffffff",
   44476 => x"ffffff",
   44477 => x"ffffff",
   44478 => x"ffffff",
   44479 => x"ffffff",
   44480 => x"ffffff",
   44481 => x"ffffff",
   44482 => x"ffffff",
   44483 => x"ffffff",
   44484 => x"ffffff",
   44485 => x"ffffff",
   44486 => x"ffffff",
   44487 => x"ffffff",
   44488 => x"ffffff",
   44489 => x"ffffff",
   44490 => x"ffffff",
   44491 => x"ffffff",
   44492 => x"ffffff",
   44493 => x"ffffff",
   44494 => x"ffffff",
   44495 => x"ffffff",
   44496 => x"ffffff",
   44497 => x"ffffff",
   44498 => x"ffffff",
   44499 => x"ffffff",
   44500 => x"ffffff",
   44501 => x"ffffff",
   44502 => x"ffffff",
   44503 => x"ffffff",
   44504 => x"ffffff",
   44505 => x"ffffeb",
   44506 => x"ad75c3",
   44507 => x"0c30c3",
   44508 => x"0c30c3",
   44509 => x"0c30c3",
   44510 => x"0c30c3",
   44511 => x"0c30c3",
   44512 => x"0c30c3",
   44513 => x"0c30c3",
   44514 => x"0c30c3",
   44515 => x"0c30c3",
   44516 => x"0c30c3",
   44517 => x"0c30c3",
   44518 => x"0c30c3",
   44519 => x"0c30c3",
   44520 => x"0c30c3",
   44521 => x"0c30c3",
   44522 => x"5d7aff",
   44523 => x"ffffff",
   44524 => x"ffffff",
   44525 => x"ffffff",
   44526 => x"ffffff",
   44527 => x"ffffff",
   44528 => x"ffffff",
   44529 => x"ffffff",
   44530 => x"ffffff",
   44531 => x"fffa80",
   44532 => x"00003f",
   44533 => x"ffffff",
   44534 => x"ffffff",
   44535 => x"ffffd5",
   44536 => x"000015",
   44537 => x"abffff",
   44538 => x"ffffff",
   44539 => x"ffffff",
   44540 => x"ffffff",
   44541 => x"ffffff",
   44542 => x"ffffff",
   44543 => x"ffffff",
   44544 => x"ffffff",
   44545 => x"ffffff",
   44546 => x"ffffff",
   44547 => x"ffffff",
   44548 => x"ffffff",
   44549 => x"fffa95",
   44550 => x"abffff",
   44551 => x"ffffff",
   44552 => x"ffffff",
   44553 => x"ffffff",
   44554 => x"ffffff",
   44555 => x"ffffff",
   44556 => x"ffffff",
   44557 => x"ffffff",
   44558 => x"ffffff",
   44559 => x"ffffff",
   44560 => x"ffffff",
   44561 => x"ffffff",
   44562 => x"ffffff",
   44563 => x"ffffff",
   44564 => x"ffffff",
   44565 => x"ffffff",
   44566 => x"ffffff",
   44567 => x"ffffff",
   44568 => x"ffffff",
   44569 => x"ffffff",
   44570 => x"ffffff",
   44571 => x"ffffff",
   44572 => x"ffffff",
   44573 => x"ffffff",
   44574 => x"ffffff",
   44575 => x"ffffff",
   44576 => x"ffffff",
   44577 => x"ffffff",
   44578 => x"ffffff",
   44579 => x"ffffff",
   44580 => x"ffffff",
   44581 => x"ffffff",
   44582 => x"ffffff",
   44583 => x"ffffff",
   44584 => x"ffffff",
   44585 => x"ffffff",
   44586 => x"ffffff",
   44587 => x"ffffff",
   44588 => x"ffffff",
   44589 => x"ffffff",
   44590 => x"ffffff",
   44591 => x"ffffff",
   44592 => x"ffffff",
   44593 => x"ffffff",
   44594 => x"ffffff",
   44595 => x"ffffff",
   44596 => x"ffffff",
   44597 => x"ffffff",
   44598 => x"ffffff",
   44599 => x"ffffff",
   44600 => x"ffffff",
   44601 => x"ffffff",
   44602 => x"ffffff",
   44603 => x"ffffff",
   44604 => x"ffffff",
   44605 => x"ffffff",
   44606 => x"ffffff",
   44607 => x"ffffff",
   44608 => x"ffffff",
   44609 => x"ffffff",
   44610 => x"ffffff",
   44611 => x"ffffff",
   44612 => x"ffffff",
   44613 => x"ffffff",
   44614 => x"ffffff",
   44615 => x"ffffff",
   44616 => x"ffffff",
   44617 => x"ffffff",
   44618 => x"ffffff",
   44619 => x"ffffff",
   44620 => x"ffffff",
   44621 => x"ffffff",
   44622 => x"ffffff",
   44623 => x"ffffff",
   44624 => x"ffffff",
   44625 => x"ffffff",
   44626 => x"ffffff",
   44627 => x"ffffff",
   44628 => x"ffffff",
   44629 => x"ffffff",
   44630 => x"ffffff",
   44631 => x"ffffff",
   44632 => x"ffffff",
   44633 => x"ffffff",
   44634 => x"ffffff",
   44635 => x"ffffff",
   44636 => x"ffffff",
   44637 => x"ffffff",
   44638 => x"ffffff",
   44639 => x"ffffff",
   44640 => x"ffffff",
   44641 => x"ffffff",
   44642 => x"ffffff",
   44643 => x"ffffff",
   44644 => x"ffffff",
   44645 => x"ffffff",
   44646 => x"ffffff",
   44647 => x"ffffff",
   44648 => x"ffffff",
   44649 => x"ffffff",
   44650 => x"ffffff",
   44651 => x"ffffff",
   44652 => x"ffffff",
   44653 => x"ffffff",
   44654 => x"ffffff",
   44655 => x"ffffff",
   44656 => x"ffffff",
   44657 => x"ffffff",
   44658 => x"ffffff",
   44659 => x"ffffff",
   44660 => x"ffffff",
   44661 => x"ffffff",
   44662 => x"ffffff",
   44663 => x"ffffff",
   44664 => x"ffffff",
   44665 => x"ffffff",
   44666 => x"fffaeb",
   44667 => x"5d70c3",
   44668 => x"0c30c3",
   44669 => x"0c30c3",
   44670 => x"0c30c3",
   44671 => x"0c30c3",
   44672 => x"0c30c3",
   44673 => x"0c30c3",
   44674 => x"0c30c3",
   44675 => x"0c30c3",
   44676 => x"0c30c3",
   44677 => x"0c30c3",
   44678 => x"0c30c3",
   44679 => x"0c30c3",
   44680 => x"0c30c3",
   44681 => x"0d75eb",
   44682 => x"ffffff",
   44683 => x"ffffff",
   44684 => x"ffffff",
   44685 => x"ffffff",
   44686 => x"ffffff",
   44687 => x"ffffff",
   44688 => x"ffffff",
   44689 => x"ffffff",
   44690 => x"ffffff",
   44691 => x"fffa80",
   44692 => x"00003f",
   44693 => x"ffffff",
   44694 => x"ffffff",
   44695 => x"fea540",
   44696 => x"000015",
   44697 => x"ffffff",
   44698 => x"ffffff",
   44699 => x"ffffff",
   44700 => x"ffffff",
   44701 => x"ffffff",
   44702 => x"ffffff",
   44703 => x"ffffff",
   44704 => x"ffffff",
   44705 => x"ffffff",
   44706 => x"ffffff",
   44707 => x"ffffff",
   44708 => x"ffffff",
   44709 => x"fffa95",
   44710 => x"abffff",
   44711 => x"ffffff",
   44712 => x"ffffff",
   44713 => x"ffffff",
   44714 => x"ffffff",
   44715 => x"ffffff",
   44716 => x"ffffff",
   44717 => x"ffffff",
   44718 => x"ffffff",
   44719 => x"ffffff",
   44720 => x"ffffff",
   44721 => x"ffffff",
   44722 => x"ffffff",
   44723 => x"ffffff",
   44724 => x"ffffff",
   44725 => x"ffffff",
   44726 => x"ffffff",
   44727 => x"ffffff",
   44728 => x"ffffff",
   44729 => x"ffffff",
   44730 => x"ffffff",
   44731 => x"ffffff",
   44732 => x"ffffff",
   44733 => x"ffffff",
   44734 => x"ffffff",
   44735 => x"ffffff",
   44736 => x"ffffff",
   44737 => x"ffffff",
   44738 => x"ffffff",
   44739 => x"ffffff",
   44740 => x"ffffff",
   44741 => x"ffffff",
   44742 => x"ffffff",
   44743 => x"ffffff",
   44744 => x"ffffff",
   44745 => x"ffffff",
   44746 => x"ffffff",
   44747 => x"ffffff",
   44748 => x"ffffff",
   44749 => x"ffffff",
   44750 => x"ffffff",
   44751 => x"ffffff",
   44752 => x"ffffff",
   44753 => x"ffffff",
   44754 => x"ffffff",
   44755 => x"ffffff",
   44756 => x"ffffff",
   44757 => x"ffffff",
   44758 => x"ffffff",
   44759 => x"ffffff",
   44760 => x"ffffff",
   44761 => x"ffffff",
   44762 => x"ffffff",
   44763 => x"ffffff",
   44764 => x"ffffff",
   44765 => x"ffffff",
   44766 => x"ffffff",
   44767 => x"ffffff",
   44768 => x"ffffff",
   44769 => x"ffffff",
   44770 => x"ffffff",
   44771 => x"ffffff",
   44772 => x"ffffff",
   44773 => x"ffffff",
   44774 => x"ffffff",
   44775 => x"ffffff",
   44776 => x"ffffff",
   44777 => x"ffffff",
   44778 => x"ffffff",
   44779 => x"ffffff",
   44780 => x"ffffff",
   44781 => x"ffffff",
   44782 => x"ffffff",
   44783 => x"ffffff",
   44784 => x"ffffff",
   44785 => x"ffffff",
   44786 => x"ffffff",
   44787 => x"ffffff",
   44788 => x"ffffff",
   44789 => x"ffffff",
   44790 => x"ffffff",
   44791 => x"ffffff",
   44792 => x"ffffff",
   44793 => x"ffffff",
   44794 => x"ffffff",
   44795 => x"ffffff",
   44796 => x"ffffff",
   44797 => x"ffffff",
   44798 => x"ffffff",
   44799 => x"ffffff",
   44800 => x"ffffff",
   44801 => x"ffffff",
   44802 => x"ffffff",
   44803 => x"ffffff",
   44804 => x"ffffff",
   44805 => x"ffffff",
   44806 => x"ffffff",
   44807 => x"ffffff",
   44808 => x"ffffff",
   44809 => x"ffffff",
   44810 => x"ffffff",
   44811 => x"ffffff",
   44812 => x"ffffff",
   44813 => x"ffffff",
   44814 => x"ffffff",
   44815 => x"ffffff",
   44816 => x"ffffff",
   44817 => x"ffffff",
   44818 => x"ffffff",
   44819 => x"ffffff",
   44820 => x"ffffff",
   44821 => x"ffffff",
   44822 => x"ffffff",
   44823 => x"ffffff",
   44824 => x"ffffff",
   44825 => x"ffffff",
   44826 => x"ffffff",
   44827 => x"febad7",
   44828 => x"5d70c3",
   44829 => x"0c30c3",
   44830 => x"0c30c3",
   44831 => x"0c30c3",
   44832 => x"0c30c3",
   44833 => x"0c30c3",
   44834 => x"0c30c3",
   44835 => x"0c30c3",
   44836 => x"0c30c3",
   44837 => x"0c30c3",
   44838 => x"0c30c3",
   44839 => x"0c30c3",
   44840 => x"0d75d7",
   44841 => x"afffff",
   44842 => x"ffffff",
   44843 => x"ffffff",
   44844 => x"ffffff",
   44845 => x"ffffff",
   44846 => x"ffffff",
   44847 => x"ffffff",
   44848 => x"ffffff",
   44849 => x"ffffff",
   44850 => x"ffffff",
   44851 => x"fffa80",
   44852 => x"00002a",
   44853 => x"aaaaaa",
   44854 => x"aaaaaa",
   44855 => x"a95000",
   44856 => x"00056a",
   44857 => x"ffffff",
   44858 => x"ffffff",
   44859 => x"ffffff",
   44860 => x"ffffff",
   44861 => x"ffffff",
   44862 => x"ffffff",
   44863 => x"ffffff",
   44864 => x"ffffff",
   44865 => x"ffffff",
   44866 => x"ffffff",
   44867 => x"ffffff",
   44868 => x"ffffff",
   44869 => x"fffa95",
   44870 => x"abffff",
   44871 => x"ffffff",
   44872 => x"ffffff",
   44873 => x"ffffff",
   44874 => x"ffffff",
   44875 => x"ffffff",
   44876 => x"ffffff",
   44877 => x"ffffff",
   44878 => x"ffffff",
   44879 => x"ffffff",
   44880 => x"ffffff",
   44881 => x"ffffff",
   44882 => x"ffffff",
   44883 => x"ffffff",
   44884 => x"ffffff",
   44885 => x"ffffff",
   44886 => x"ffffff",
   44887 => x"ffffff",
   44888 => x"ffffff",
   44889 => x"ffffff",
   44890 => x"ffffff",
   44891 => x"ffffff",
   44892 => x"ffffff",
   44893 => x"ffffff",
   44894 => x"ffffff",
   44895 => x"ffffff",
   44896 => x"ffffff",
   44897 => x"ffffff",
   44898 => x"ffffff",
   44899 => x"ffffff",
   44900 => x"ffffff",
   44901 => x"ffffff",
   44902 => x"ffffff",
   44903 => x"ffffff",
   44904 => x"ffffff",
   44905 => x"ffffff",
   44906 => x"ffffff",
   44907 => x"ffffff",
   44908 => x"ffffff",
   44909 => x"ffffff",
   44910 => x"ffffff",
   44911 => x"ffffff",
   44912 => x"ffffff",
   44913 => x"ffffff",
   44914 => x"ffffff",
   44915 => x"ffffff",
   44916 => x"ffffff",
   44917 => x"ffffff",
   44918 => x"ffffff",
   44919 => x"ffffff",
   44920 => x"ffffff",
   44921 => x"ffffff",
   44922 => x"ffffff",
   44923 => x"ffffff",
   44924 => x"ffffff",
   44925 => x"ffffff",
   44926 => x"ffffff",
   44927 => x"ffffff",
   44928 => x"ffffff",
   44929 => x"ffffff",
   44930 => x"ffffff",
   44931 => x"ffffff",
   44932 => x"ffffff",
   44933 => x"ffffff",
   44934 => x"ffffff",
   44935 => x"ffffff",
   44936 => x"ffffff",
   44937 => x"ffffff",
   44938 => x"ffffff",
   44939 => x"ffffff",
   44940 => x"ffffff",
   44941 => x"ffffff",
   44942 => x"ffffff",
   44943 => x"ffffff",
   44944 => x"ffffff",
   44945 => x"ffffff",
   44946 => x"ffffff",
   44947 => x"ffffff",
   44948 => x"ffffff",
   44949 => x"ffffff",
   44950 => x"ffffff",
   44951 => x"ffffff",
   44952 => x"ffffff",
   44953 => x"ffffff",
   44954 => x"ffffff",
   44955 => x"ffffff",
   44956 => x"ffffff",
   44957 => x"ffffff",
   44958 => x"ffffff",
   44959 => x"ffffff",
   44960 => x"ffffff",
   44961 => x"ffffff",
   44962 => x"ffffff",
   44963 => x"ffffff",
   44964 => x"ffffff",
   44965 => x"ffffff",
   44966 => x"ffffff",
   44967 => x"ffffff",
   44968 => x"ffffff",
   44969 => x"ffffff",
   44970 => x"ffffff",
   44971 => x"ffffff",
   44972 => x"ffffff",
   44973 => x"ffffff",
   44974 => x"ffffff",
   44975 => x"ffffff",
   44976 => x"ffffff",
   44977 => x"ffffff",
   44978 => x"ffffff",
   44979 => x"ffffff",
   44980 => x"ffffff",
   44981 => x"ffffff",
   44982 => x"ffffff",
   44983 => x"ffffff",
   44984 => x"ffffff",
   44985 => x"ffffff",
   44986 => x"ffffff",
   44987 => x"ffffff",
   44988 => x"febad7",
   44989 => x"5c30c3",
   44990 => x"0c30c3",
   44991 => x"0c30c3",
   44992 => x"0c30c3",
   44993 => x"0c30c3",
   44994 => x"0c30c3",
   44995 => x"0c30c3",
   44996 => x"0c30c3",
   44997 => x"0c30c3",
   44998 => x"0c30c3",
   44999 => x"0d75d7",
   45000 => x"aebfff",
   45001 => x"ffffff",
   45002 => x"ffffff",
   45003 => x"ffffff",
   45004 => x"ffffff",
   45005 => x"ffffff",
   45006 => x"ffffff",
   45007 => x"ffffff",
   45008 => x"ffffff",
   45009 => x"ffffff",
   45010 => x"ffffff",
   45011 => x"fffa80",
   45012 => x"000000",
   45013 => x"000000",
   45014 => x"000000",
   45015 => x"000000",
   45016 => x"000abf",
   45017 => x"ffffff",
   45018 => x"ffffff",
   45019 => x"ffffff",
   45020 => x"ffffff",
   45021 => x"ffffff",
   45022 => x"ffffff",
   45023 => x"ffffff",
   45024 => x"ffffff",
   45025 => x"ffffff",
   45026 => x"ffffff",
   45027 => x"ffffff",
   45028 => x"ffffff",
   45029 => x"fffa95",
   45030 => x"abffff",
   45031 => x"ffffff",
   45032 => x"ffffff",
   45033 => x"ffffff",
   45034 => x"ffffff",
   45035 => x"ffffff",
   45036 => x"ffffff",
   45037 => x"ffffff",
   45038 => x"ffffff",
   45039 => x"ffffff",
   45040 => x"ffffff",
   45041 => x"ffffff",
   45042 => x"ffffff",
   45043 => x"ffffff",
   45044 => x"ffffff",
   45045 => x"ffffff",
   45046 => x"ffffff",
   45047 => x"ffffff",
   45048 => x"ffffff",
   45049 => x"ffffff",
   45050 => x"ffffff",
   45051 => x"ffffff",
   45052 => x"ffffff",
   45053 => x"ffffff",
   45054 => x"ffffff",
   45055 => x"ffffff",
   45056 => x"ffffff",
   45057 => x"ffffff",
   45058 => x"ffffff",
   45059 => x"ffffff",
   45060 => x"ffffff",
   45061 => x"ffffff",
   45062 => x"ffffff",
   45063 => x"ffffff",
   45064 => x"ffffff",
   45065 => x"ffffff",
   45066 => x"ffffff",
   45067 => x"ffffff",
   45068 => x"ffffff",
   45069 => x"ffffff",
   45070 => x"ffffff",
   45071 => x"ffffff",
   45072 => x"ffffff",
   45073 => x"ffffff",
   45074 => x"ffffff",
   45075 => x"ffffff",
   45076 => x"ffffff",
   45077 => x"ffffff",
   45078 => x"ffffff",
   45079 => x"ffffff",
   45080 => x"ffffff",
   45081 => x"ffffff",
   45082 => x"ffffff",
   45083 => x"ffffff",
   45084 => x"ffffff",
   45085 => x"ffffff",
   45086 => x"ffffff",
   45087 => x"ffffff",
   45088 => x"ffffff",
   45089 => x"ffffff",
   45090 => x"ffffff",
   45091 => x"ffffff",
   45092 => x"ffffff",
   45093 => x"ffffff",
   45094 => x"ffffff",
   45095 => x"ffffff",
   45096 => x"ffffff",
   45097 => x"ffffff",
   45098 => x"ffffff",
   45099 => x"ffffff",
   45100 => x"ffffff",
   45101 => x"ffffff",
   45102 => x"ffffff",
   45103 => x"ffffff",
   45104 => x"ffffff",
   45105 => x"ffffff",
   45106 => x"ffffff",
   45107 => x"ffffff",
   45108 => x"ffffff",
   45109 => x"ffffff",
   45110 => x"ffffff",
   45111 => x"ffffff",
   45112 => x"ffffff",
   45113 => x"ffffff",
   45114 => x"ffffff",
   45115 => x"ffffff",
   45116 => x"ffffff",
   45117 => x"ffffff",
   45118 => x"ffffff",
   45119 => x"ffffff",
   45120 => x"ffffff",
   45121 => x"ffffff",
   45122 => x"ffffff",
   45123 => x"ffffff",
   45124 => x"ffffff",
   45125 => x"ffffff",
   45126 => x"ffffff",
   45127 => x"ffffff",
   45128 => x"ffffff",
   45129 => x"ffffff",
   45130 => x"ffffff",
   45131 => x"ffffff",
   45132 => x"ffffff",
   45133 => x"ffffff",
   45134 => x"ffffff",
   45135 => x"ffffff",
   45136 => x"ffffff",
   45137 => x"ffffff",
   45138 => x"ffffff",
   45139 => x"ffffff",
   45140 => x"ffffff",
   45141 => x"ffffff",
   45142 => x"ffffff",
   45143 => x"ffffff",
   45144 => x"ffffff",
   45145 => x"ffffff",
   45146 => x"ffffff",
   45147 => x"ffffff",
   45148 => x"ffffff",
   45149 => x"febad7",
   45150 => x"5d75c3",
   45151 => x"0c30c3",
   45152 => x"0c30c3",
   45153 => x"0c30c3",
   45154 => x"0c30c3",
   45155 => x"0c30c3",
   45156 => x"0c30c3",
   45157 => x"0c30c3",
   45158 => x"5d75d7",
   45159 => x"aebfff",
   45160 => x"ffffff",
   45161 => x"ffffff",
   45162 => x"ffffff",
   45163 => x"ffffff",
   45164 => x"ffffff",
   45165 => x"ffffff",
   45166 => x"ffffff",
   45167 => x"ffffff",
   45168 => x"ffffff",
   45169 => x"ffffff",
   45170 => x"ffffff",
   45171 => x"fffa80",
   45172 => x"000000",
   45173 => x"000000",
   45174 => x"000000",
   45175 => x"000000",
   45176 => x"56afff",
   45177 => x"ffffff",
   45178 => x"ffffff",
   45179 => x"ffffff",
   45180 => x"ffffff",
   45181 => x"ffffff",
   45182 => x"ffffff",
   45183 => x"ffffff",
   45184 => x"ffffff",
   45185 => x"ffffff",
   45186 => x"ffffff",
   45187 => x"ffffff",
   45188 => x"ffffff",
   45189 => x"fffa95",
   45190 => x"abffff",
   45191 => x"ffffff",
   45192 => x"ffffff",
   45193 => x"ffffff",
   45194 => x"ffffff",
   45195 => x"ffffff",
   45196 => x"ffffff",
   45197 => x"ffffff",
   45198 => x"ffffff",
   45199 => x"ffffff",
   45200 => x"ffffff",
   45201 => x"ffffff",
   45202 => x"ffffff",
   45203 => x"ffffff",
   45204 => x"ffffff",
   45205 => x"ffffff",
   45206 => x"ffffff",
   45207 => x"ffffff",
   45208 => x"ffffff",
   45209 => x"ffffff",
   45210 => x"ffffff",
   45211 => x"ffffff",
   45212 => x"ffffff",
   45213 => x"ffffff",
   45214 => x"ffffff",
   45215 => x"ffffff",
   45216 => x"ffffff",
   45217 => x"ffffff",
   45218 => x"ffffff",
   45219 => x"ffffff",
   45220 => x"ffffff",
   45221 => x"ffffff",
   45222 => x"ffffff",
   45223 => x"ffffff",
   45224 => x"ffffff",
   45225 => x"ffffff",
   45226 => x"ffffff",
   45227 => x"ffffff",
   45228 => x"ffffff",
   45229 => x"ffffff",
   45230 => x"ffffff",
   45231 => x"ffffff",
   45232 => x"ffffff",
   45233 => x"ffffff",
   45234 => x"ffffff",
   45235 => x"ffffff",
   45236 => x"ffffff",
   45237 => x"ffffff",
   45238 => x"ffffff",
   45239 => x"ffffff",
   45240 => x"ffffff",
   45241 => x"ffffff",
   45242 => x"ffffff",
   45243 => x"ffffff",
   45244 => x"ffffff",
   45245 => x"ffffff",
   45246 => x"ffffff",
   45247 => x"ffffff",
   45248 => x"ffffff",
   45249 => x"ffffff",
   45250 => x"ffffff",
   45251 => x"ffffff",
   45252 => x"ffffff",
   45253 => x"ffffff",
   45254 => x"ffffff",
   45255 => x"ffffff",
   45256 => x"ffffff",
   45257 => x"ffffff",
   45258 => x"ffffff",
   45259 => x"ffffff",
   45260 => x"ffffff",
   45261 => x"ffffff",
   45262 => x"ffffff",
   45263 => x"ffffff",
   45264 => x"ffffff",
   45265 => x"ffffff",
   45266 => x"ffffff",
   45267 => x"ffffff",
   45268 => x"ffffff",
   45269 => x"ffffff",
   45270 => x"ffffff",
   45271 => x"ffffff",
   45272 => x"ffffff",
   45273 => x"ffffff",
   45274 => x"ffffff",
   45275 => x"ffffff",
   45276 => x"ffffff",
   45277 => x"ffffff",
   45278 => x"ffffff",
   45279 => x"ffffff",
   45280 => x"ffffff",
   45281 => x"ffffff",
   45282 => x"ffffff",
   45283 => x"ffffff",
   45284 => x"ffffff",
   45285 => x"ffffff",
   45286 => x"ffffff",
   45287 => x"ffffff",
   45288 => x"ffffff",
   45289 => x"ffffff",
   45290 => x"ffffff",
   45291 => x"ffffff",
   45292 => x"ffffff",
   45293 => x"ffffff",
   45294 => x"ffffff",
   45295 => x"ffffff",
   45296 => x"ffffff",
   45297 => x"ffffff",
   45298 => x"ffffff",
   45299 => x"ffffff",
   45300 => x"ffffff",
   45301 => x"ffffff",
   45302 => x"ffffff",
   45303 => x"ffffff",
   45304 => x"ffffff",
   45305 => x"ffffff",
   45306 => x"ffffff",
   45307 => x"ffffff",
   45308 => x"ffffff",
   45309 => x"ffffff",
   45310 => x"fffaeb",
   45311 => x"ad75d7",
   45312 => x"5d70c3",
   45313 => x"0c30c3",
   45314 => x"0c30c3",
   45315 => x"0c30c3",
   45316 => x"0d75d7",
   45317 => x"5d7aeb",
   45318 => x"afffff",
   45319 => x"ffffff",
   45320 => x"ffffff",
   45321 => x"ffffff",
   45322 => x"ffffff",
   45323 => x"ffffff",
   45324 => x"ffffff",
   45325 => x"ffffff",
   45326 => x"ffffff",
   45327 => x"ffffff",
   45328 => x"ffffff",
   45329 => x"ffffff",
   45330 => x"ffffff",
   45331 => x"fffa95",
   45332 => x"000000",
   45333 => x"000000",
   45334 => x"000000",
   45335 => x"01556a",
   45336 => x"ffffff",
   45337 => x"ffffff",
   45338 => x"ffffff",
   45339 => x"ffffff",
   45340 => x"ffffff",
   45341 => x"ffffff",
   45342 => x"ffffff",
   45343 => x"ffffff",
   45344 => x"ffffff",
   45345 => x"ffffff",
   45346 => x"ffffff",
   45347 => x"ffffff",
   45348 => x"ffffff",
   45349 => x"fffa95",
   45350 => x"abffff",
   45351 => x"ffffff",
   45352 => x"ffffff",
   45353 => x"ffffff",
   45354 => x"ffffff",
   45355 => x"ffffff",
   45356 => x"ffffff",
   45357 => x"ffffff",
   45358 => x"ffffff",
   45359 => x"ffffff",
   45360 => x"ffffff",
   45361 => x"ffffff",
   45362 => x"ffffff",
   45363 => x"ffffff",
   45364 => x"ffffff",
   45365 => x"ffffff",
   45366 => x"ffffff",
   45367 => x"ffffff",
   45368 => x"ffffff",
   45369 => x"ffffff",
   45370 => x"ffffff",
   45371 => x"ffffff",
   45372 => x"ffffff",
   45373 => x"ffffff",
   45374 => x"ffffff",
   45375 => x"ffffff",
   45376 => x"ffffff",
   45377 => x"ffffff",
   45378 => x"ffffff",
   45379 => x"ffffff",
   45380 => x"ffffff",
   45381 => x"ffffff",
   45382 => x"ffffff",
   45383 => x"ffffff",
   45384 => x"ffffff",
   45385 => x"ffffff",
   45386 => x"ffffff",
   45387 => x"ffffff",
   45388 => x"ffffff",
   45389 => x"ffffff",
   45390 => x"ffffff",
   45391 => x"ffffff",
   45392 => x"ffffff",
   45393 => x"ffffff",
   45394 => x"ffffff",
   45395 => x"ffffff",
   45396 => x"ffffff",
   45397 => x"ffffff",
   45398 => x"ffffff",
   45399 => x"ffffff",
   45400 => x"ffffff",
   45401 => x"ffffff",
   45402 => x"ffffff",
   45403 => x"ffffff",
   45404 => x"ffffff",
   45405 => x"ffffff",
   45406 => x"ffffff",
   45407 => x"ffffff",
   45408 => x"ffffff",
   45409 => x"ffffff",
   45410 => x"ffffff",
   45411 => x"ffffff",
   45412 => x"ffffff",
   45413 => x"ffffff",
   45414 => x"ffffff",
   45415 => x"ffffff",
   45416 => x"ffffff",
   45417 => x"ffffff",
   45418 => x"ffffff",
   45419 => x"ffffff",
   45420 => x"ffffff",
   45421 => x"ffffff",
   45422 => x"ffffff",
   45423 => x"ffffff",
   45424 => x"ffffff",
   45425 => x"ffffff",
   45426 => x"ffffff",
   45427 => x"ffffff",
   45428 => x"ffffff",
   45429 => x"ffffff",
   45430 => x"ffffff",
   45431 => x"ffffff",
   45432 => x"ffffff",
   45433 => x"ffffff",
   45434 => x"ffffff",
   45435 => x"ffffff",
   45436 => x"ffffff",
   45437 => x"ffffff",
   45438 => x"ffffff",
   45439 => x"ffffff",
   45440 => x"ffffff",
   45441 => x"ffffff",
   45442 => x"ffffff",
   45443 => x"ffffff",
   45444 => x"ffffff",
   45445 => x"ffffff",
   45446 => x"ffffff",
   45447 => x"ffffff",
   45448 => x"ffffff",
   45449 => x"ffffff",
   45450 => x"ffffff",
   45451 => x"ffffff",
   45452 => x"ffffff",
   45453 => x"ffffff",
   45454 => x"ffffff",
   45455 => x"ffffff",
   45456 => x"ffffff",
   45457 => x"ffffff",
   45458 => x"ffffff",
   45459 => x"ffffff",
   45460 => x"ffffff",
   45461 => x"ffffff",
   45462 => x"ffffff",
   45463 => x"ffffff",
   45464 => x"ffffff",
   45465 => x"ffffff",
   45466 => x"ffffff",
   45467 => x"ffffff",
   45468 => x"ffffff",
   45469 => x"ffffff",
   45470 => x"ffffff",
   45471 => x"ffffff",
   45472 => x"fffaeb",
   45473 => x"aebaeb",
   45474 => x"aebaeb",
   45475 => x"aebaeb",
   45476 => x"ffffff",
   45477 => x"ffffff",
   45478 => x"ffffff",
   45479 => x"ffffff",
   45480 => x"ffffff",
   45481 => x"ffffff",
   45482 => x"ffffff",
   45483 => x"ffffff",
   45484 => x"ffffff",
   45485 => x"ffffff",
   45486 => x"ffffff",
   45487 => x"ffffff",
   45488 => x"ffffff",
   45489 => x"ffffff",
   45490 => x"ffffff",
   45491 => x"ffffea",
   45492 => x"aaaaaa",
   45493 => x"aaaaaa",
   45494 => x"aaaaaa",
   45495 => x"abffff",
   45496 => x"ffffff",
   45497 => x"ffffff",
   45498 => x"ffffff",
   45499 => x"ffffff",
   45500 => x"ffffff",
   45501 => x"ffffff",
   45502 => x"ffffff",
   45503 => x"ffffff",
   45504 => x"ffffff",
   45505 => x"ffffff",
   45506 => x"ffffff",
   45507 => x"ffffff",
   45508 => x"ffffff",
   45509 => x"fffa95",
   45510 => x"abffff",
   45511 => x"ffffff",
   45512 => x"ffffff",
   45513 => x"ffffff",
   45514 => x"ffffff",
   45515 => x"ffffff",
   45516 => x"ffffff",
   45517 => x"ffffff",
   45518 => x"ffffff",
   45519 => x"ffffff",
   45520 => x"ffffff",
   45521 => x"ffffff",
   45522 => x"ffffff",
   45523 => x"ffffff",
   45524 => x"ffffff",
   45525 => x"ffffff",
   45526 => x"ffffff",
   45527 => x"ffffff",
   45528 => x"ffffff",
   45529 => x"ffffff",
   45530 => x"ffffff",
   45531 => x"ffffff",
   45532 => x"ffffff",
   45533 => x"ffffff",
   45534 => x"ffffff",
   45535 => x"ffffff",
   45536 => x"ffffff",
   45537 => x"ffffff",
   45538 => x"ffffff",
   45539 => x"ffffff",
   45540 => x"ffffff",
   45541 => x"ffffff",
   45542 => x"ffffff",
   45543 => x"ffffff",
   45544 => x"ffffff",
   45545 => x"ffffff",
   45546 => x"ffffff",
   45547 => x"ffffff",
   45548 => x"ffffff",
   45549 => x"ffffff",
   45550 => x"ffffff",
   45551 => x"ffffff",
   45552 => x"ffffff",
   45553 => x"ffffff",
   45554 => x"ffffff",
   45555 => x"ffffff",
   45556 => x"ffffff",
   45557 => x"ffffff",
   45558 => x"ffffff",
   45559 => x"ffffff",
   45560 => x"ffffff",
   45561 => x"ffffff",
   45562 => x"ffffff",
   45563 => x"ffffff",
   45564 => x"ffffff",
   45565 => x"ffffff",
   45566 => x"ffffff",
   45567 => x"ffffff",
   45568 => x"ffffff",
   45569 => x"ffffff",
   45570 => x"ffffff",
   45571 => x"ffffff",
   45572 => x"ffffff",
   45573 => x"ffffff",
   45574 => x"ffffff",
   45575 => x"ffffff",
   45576 => x"ffffff",
   45577 => x"ffffff",
   45578 => x"ffffff",
   45579 => x"ffffff",
   45580 => x"ffffff",
   45581 => x"ffffff",
   45582 => x"ffffff",
   45583 => x"ffffff",
   45584 => x"ffffff",
   45585 => x"ffffff",
   45586 => x"ffffff",
   45587 => x"ffffff",
   45588 => x"ffffff",
   45589 => x"ffffff",
   45590 => x"ffffff",
   45591 => x"ffffff",
   45592 => x"ffffff",
   45593 => x"ffffff",
   45594 => x"ffffff",
   45595 => x"ffffff",
   45596 => x"ffffff",
   45597 => x"ffffff",
   45598 => x"ffffff",
   45599 => x"ffffff",
   45600 => x"ffffff",
   45601 => x"ffffff",
   45602 => x"ffffff",
   45603 => x"ffffff",
   45604 => x"ffffff",
   45605 => x"ffffff",
   45606 => x"ffffff",
   45607 => x"ffffff",
   45608 => x"ffffff",
   45609 => x"ffffff",
   45610 => x"ffffff",
   45611 => x"ffffff",
   45612 => x"ffffff",
   45613 => x"ffffff",
   45614 => x"ffffff",
   45615 => x"ffffff",
   45616 => x"ffffff",
   45617 => x"ffffff",
   45618 => x"ffffff",
   45619 => x"ffffff",
   45620 => x"ffffff",
   45621 => x"ffffff",
   45622 => x"ffffff",
   45623 => x"ffffff",
   45624 => x"ffffff",
   45625 => x"ffffff",
   45626 => x"ffffff",
   45627 => x"ffffff",
   45628 => x"ffffff",
   45629 => x"ffffff",
   45630 => x"ffffff",
   45631 => x"ffffff",
   45632 => x"ffffff",
   45633 => x"ffffff",
   45634 => x"ffffff",
   45635 => x"ffffff",
   45636 => x"ffffff",
   45637 => x"ffffff",
   45638 => x"ffffff",
   45639 => x"ffffff",
   45640 => x"ffffff",
   45641 => x"ffffff",
   45642 => x"ffffff",
   45643 => x"ffffff",
   45644 => x"ffffff",
   45645 => x"ffffff",
   45646 => x"ffffff",
   45647 => x"ffffff",
   45648 => x"ffffff",
   45649 => x"ffffff",
   45650 => x"ffffff",
   45651 => x"ffffff",
   45652 => x"ffffff",
   45653 => x"ffffff",
   45654 => x"ffffff",
   45655 => x"ffffff",
   45656 => x"ffffff",
   45657 => x"ffffff",
   45658 => x"ffffff",
   45659 => x"ffffff",
   45660 => x"ffffff",
   45661 => x"ffffff",
   45662 => x"ffffff",
   45663 => x"ffffff",
   45664 => x"ffffff",
   45665 => x"ffffff",
   45666 => x"ffffff",
   45667 => x"ffffff",
   45668 => x"ffffff",
   45669 => x"fffa95",
   45670 => x"abffff",
   45671 => x"ffffff",
   45672 => x"ffffff",
   45673 => x"ffffff",
   45674 => x"ffffff",
   45675 => x"ffffff",
   45676 => x"ffffff",
   45677 => x"ffffff",
   45678 => x"ffffff",
   45679 => x"ffffff",
   45680 => x"ffffff",
   45681 => x"ffffff",
   45682 => x"ffffff",
   45683 => x"ffffff",
   45684 => x"ffffff",
   45685 => x"ffffff",
   45686 => x"ffffff",
   45687 => x"ffffff",
   45688 => x"ffffff",
   45689 => x"ffffff",
   45690 => x"ffffff",
   45691 => x"ffffff",
   45692 => x"ffffff",
   45693 => x"ffffff",
   45694 => x"ffffff",
   45695 => x"ffffff",
   45696 => x"ffffff",
   45697 => x"ffffff",
   45698 => x"ffffff",
   45699 => x"ffffff",
   45700 => x"ffffff",
   45701 => x"ffffff",
   45702 => x"ffffff",
   45703 => x"ffffff",
   45704 => x"ffffff",
   45705 => x"ffffff",
   45706 => x"ffffff",
   45707 => x"ffffff",
   45708 => x"ffffff",
   45709 => x"ffffff",
   45710 => x"ffffff",
   45711 => x"ffffff",
   45712 => x"ffffff",
   45713 => x"ffffff",
   45714 => x"ffffff",
   45715 => x"ffffff",
   45716 => x"ffffff",
   45717 => x"ffffff",
   45718 => x"ffffff",
   45719 => x"ffffff",
   45720 => x"ffffff",
   45721 => x"ffffff",
   45722 => x"ffffff",
   45723 => x"ffffff",
   45724 => x"ffffff",
   45725 => x"ffffff",
   45726 => x"ffffff",
   45727 => x"ffffff",
   45728 => x"ffffff",
   45729 => x"ffffff",
   45730 => x"ffffff",
   45731 => x"ffffff",
   45732 => x"ffffff",
   45733 => x"ffffff",
   45734 => x"ffffff",
   45735 => x"ffffff",
   45736 => x"ffffff",
   45737 => x"ffffff",
   45738 => x"ffffff",
   45739 => x"ffffff",
   45740 => x"ffffff",
   45741 => x"ffffff",
   45742 => x"ffffff",
   45743 => x"ffffff",
   45744 => x"ffffff",
   45745 => x"ffffff",
   45746 => x"ffffff",
   45747 => x"ffffff",
   45748 => x"ffffff",
   45749 => x"ffffff",
   45750 => x"ffffff",
   45751 => x"ffffff",
   45752 => x"ffffff",
   45753 => x"ffffff",
   45754 => x"ffffff",
   45755 => x"ffffff",
   45756 => x"ffffff",
   45757 => x"ffffff",
   45758 => x"ffffff",
   45759 => x"ffffff",
   45760 => x"ffffff",
   45761 => x"ffffff",
   45762 => x"ffffff",
   45763 => x"ffffff",
   45764 => x"ffffff",
   45765 => x"ffffff",
   45766 => x"ffffff",
   45767 => x"ffffff",
   45768 => x"ffffff",
   45769 => x"ffffff",
   45770 => x"ffffff",
   45771 => x"ffffff",
   45772 => x"ffffff",
   45773 => x"ffffff",
   45774 => x"ffffff",
   45775 => x"ffffff",
   45776 => x"ffffff",
   45777 => x"ffffff",
   45778 => x"ffffff",
   45779 => x"ffffff",
   45780 => x"ffffff",
   45781 => x"ffffff",
   45782 => x"ffffff",
   45783 => x"ffffff",
   45784 => x"ffffff",
   45785 => x"ffffff",
   45786 => x"ffffff",
   45787 => x"ffffff",
   45788 => x"ffffff",
   45789 => x"ffffff",
   45790 => x"ffffff",
   45791 => x"ffffff",
   45792 => x"ffffff",
   45793 => x"ffffff",
   45794 => x"ffffff",
   45795 => x"ffffff",
   45796 => x"ffffff",
   45797 => x"ffffff",
   45798 => x"ffffff",
   45799 => x"ffffff",
   45800 => x"ffffff",
   45801 => x"ffffff",
   45802 => x"ffffff",
   45803 => x"ffffff",
   45804 => x"ffffff",
   45805 => x"ffffff",
   45806 => x"ffffff",
   45807 => x"ffffff",
   45808 => x"ffffff",
   45809 => x"ffffff",
   45810 => x"ffffff",
   45811 => x"ffffff",
   45812 => x"ffffff",
   45813 => x"ffffff",
   45814 => x"ffffff",
   45815 => x"ffffff",
   45816 => x"ffffff",
   45817 => x"ffffff",
   45818 => x"ffffff",
   45819 => x"ffffff",
   45820 => x"ffffff",
   45821 => x"ffffff",
   45822 => x"ffffff",
   45823 => x"ffffff",
   45824 => x"ffffff",
   45825 => x"ffffff",
   45826 => x"ffffff",
   45827 => x"ffffff",
   45828 => x"ffffff",
   45829 => x"fffa95",
   45830 => x"abffff",
   45831 => x"ffffff",
   45832 => x"ffffff",
   45833 => x"ffffff",
   45834 => x"ffffff",
   45835 => x"ffffff",
   45836 => x"ffffff",
   45837 => x"ffffff",
   45838 => x"ffffff",
   45839 => x"ffffff",
   45840 => x"ffffff",
   45841 => x"ffffff",
   45842 => x"ffffff",
   45843 => x"ffffff",
   45844 => x"ffffff",
   45845 => x"ffffff",
   45846 => x"ffffff",
   45847 => x"ffffff",
   45848 => x"ffffff",
   45849 => x"ffffff",
   45850 => x"ffffff",
   45851 => x"ffffff",
   45852 => x"ffffff",
   45853 => x"ffffff",
   45854 => x"ffffff",
   45855 => x"ffffff",
   45856 => x"ffffff",
   45857 => x"ffffff",
   45858 => x"ffffff",
   45859 => x"ffffff",
   45860 => x"ffffff",
   45861 => x"ffffff",
   45862 => x"ffffff",
   45863 => x"ffffff",
   45864 => x"ffffff",
   45865 => x"ffffff",
   45866 => x"ffffff",
   45867 => x"ffffff",
   45868 => x"ffffff",
   45869 => x"ffffff",
   45870 => x"ffffff",
   45871 => x"ffffff",
   45872 => x"ffffff",
   45873 => x"ffffff",
   45874 => x"ffffff",
   45875 => x"ffffff",
   45876 => x"ffffff",
   45877 => x"ffffff",
   45878 => x"ffffff",
   45879 => x"ffffff",
   45880 => x"ffffff",
   45881 => x"ffffff",
   45882 => x"ffffff",
   45883 => x"ffffff",
   45884 => x"ffffff",
   45885 => x"ffffff",
   45886 => x"ffffff",
   45887 => x"ffffff",
   45888 => x"ffffff",
   45889 => x"ffffff",
   45890 => x"ffffff",
   45891 => x"ffffff",
   45892 => x"ffffff",
   45893 => x"ffffff",
   45894 => x"ffffff",
   45895 => x"ffffff",
   45896 => x"ffffff",
   45897 => x"ffffff",
   45898 => x"ffffff",
   45899 => x"ffffff",
   45900 => x"ffffff",
   45901 => x"ffffff",
   45902 => x"ffffff",
   45903 => x"ffffff",
   45904 => x"ffffff",
   45905 => x"ffffff",
   45906 => x"ffffff",
   45907 => x"ffffff",
   45908 => x"ffffff",
   45909 => x"ffffff",
   45910 => x"ffffff",
   45911 => x"ffffff",
   45912 => x"ffffff",
   45913 => x"ffffff",
   45914 => x"ffffff",
   45915 => x"ffffff",
   45916 => x"ffffff",
   45917 => x"ffffff",
   45918 => x"ffffff",
   45919 => x"ffffff",
   45920 => x"ffffff",
   45921 => x"ffffff",
   45922 => x"ffffff",
   45923 => x"ffffff",
   45924 => x"ffffff",
   45925 => x"ffffff",
   45926 => x"ffffff",
   45927 => x"ffffff",
   45928 => x"ffffff",
   45929 => x"ffffff",
   45930 => x"ffffff",
   45931 => x"ffffff",
   45932 => x"ffffff",
   45933 => x"ffffff",
   45934 => x"ffffff",
   45935 => x"ffffff",
   45936 => x"ffffff",
   45937 => x"ffffff",
   45938 => x"ffffff",
   45939 => x"ffffff",
   45940 => x"ffffff",
   45941 => x"ffffff",
   45942 => x"ffffff",
   45943 => x"ffffff",
   45944 => x"ffffff",
   45945 => x"ffffff",
   45946 => x"ffffff",
   45947 => x"ffffff",
   45948 => x"ffffff",
   45949 => x"ffffff",
   45950 => x"ffffff",
   45951 => x"ffffff",
   45952 => x"ffffff",
   45953 => x"ffffff",
   45954 => x"ffffff",
   45955 => x"ffffff",
   45956 => x"ffffff",
   45957 => x"ffffff",
   45958 => x"ffffff",
   45959 => x"ffffff",
   45960 => x"ffffff",
   45961 => x"ffffff",
   45962 => x"ffffff",
   45963 => x"ffffff",
   45964 => x"ffffff",
   45965 => x"ffffff",
   45966 => x"ffffff",
   45967 => x"ffffff",
   45968 => x"ffffff",
   45969 => x"ffffff",
   45970 => x"ffffff",
   45971 => x"ffffff",
   45972 => x"ffffff",
   45973 => x"ffffff",
   45974 => x"ffffff",
   45975 => x"ffffff",
   45976 => x"ffffff",
   45977 => x"ffffff",
   45978 => x"ffffff",
   45979 => x"ffffff",
   45980 => x"ffffff",
   45981 => x"ffffff",
   45982 => x"ffffff",
   45983 => x"ffffff",
   45984 => x"ffffff",
   45985 => x"ffffff",
   45986 => x"ffffff",
   45987 => x"ffffff",
   45988 => x"ffffff",
   45989 => x"fffa95",
   45990 => x"abffff",
   45991 => x"ffffff",
   45992 => x"ffffff",
   45993 => x"ffffff",
   45994 => x"ffffff",
   45995 => x"ffffff",
   45996 => x"ffffff",
   45997 => x"ffffff",
   45998 => x"ffffff",
   45999 => x"ffffff",
   46000 => x"ffffff",
   46001 => x"ffffff",
   46002 => x"ffffff",
   46003 => x"ffffff",
   46004 => x"ffffff",
   46005 => x"ffffff",
   46006 => x"ffffff",
   46007 => x"ffffff",
   46008 => x"ffffff",
   46009 => x"ffffff",
   46010 => x"ffffff",
   46011 => x"ffffff",
   46012 => x"ffffff",
   46013 => x"ffffff",
   46014 => x"ffffff",
   46015 => x"ffffff",
   46016 => x"ffffff",
   46017 => x"ffffff",
   46018 => x"ffffff",
   46019 => x"ffffff",
   46020 => x"ffffff",
   46021 => x"ffffff",
   46022 => x"ffffff",
   46023 => x"ffffff",
   46024 => x"ffffff",
   46025 => x"ffffff",
   46026 => x"ffffff",
   46027 => x"ffffff",
   46028 => x"ffffff",
   46029 => x"ffffff",
   46030 => x"ffffff",
   46031 => x"ffffff",
   46032 => x"ffffff",
   46033 => x"ffffff",
   46034 => x"ffffff",
   46035 => x"ffffff",
   46036 => x"ffffff",
   46037 => x"ffffff",
   46038 => x"ffffff",
   46039 => x"ffffff",
   46040 => x"ffffff",
   46041 => x"ffffff",
   46042 => x"ffffff",
   46043 => x"ffffff",
   46044 => x"ffffff",
   46045 => x"ffffff",
   46046 => x"ffffff",
   46047 => x"ffffff",
   46048 => x"ffffff",
   46049 => x"ffffff",
   46050 => x"ffffff",
   46051 => x"ffffff",
   46052 => x"ffffff",
   46053 => x"ffffff",
   46054 => x"ffffff",
   46055 => x"ffffff",
   46056 => x"ffffff",
   46057 => x"ffffff",
   46058 => x"ffffff",
   46059 => x"ffffff",
   46060 => x"ffffff",
   46061 => x"ffffff",
   46062 => x"ffffff",
   46063 => x"ffffff",
   46064 => x"ffffff",
   46065 => x"ffffff",
   46066 => x"ffffff",
   46067 => x"ffffff",
   46068 => x"ffffff",
   46069 => x"ffffff",
   46070 => x"ffffff",
   46071 => x"ffffff",
   46072 => x"ffffff",
   46073 => x"ffffff",
   46074 => x"ffffff",
   46075 => x"ffffff",
   46076 => x"ffffff",
   46077 => x"ffffff",
   46078 => x"ffffff",
   46079 => x"ffffff",
   46080 => x"ffffff",
   46081 => x"ffffff",
   46082 => x"ffffff",
   46083 => x"ffffff",
   46084 => x"ffffff",
   46085 => x"ffffff",
   46086 => x"ffffff",
   46087 => x"ffffff",
   46088 => x"ffffff",
   46089 => x"ffffff",
   46090 => x"ffffff",
   46091 => x"ffffff",
   46092 => x"ffffff",
   46093 => x"ffffff",
   46094 => x"ffffff",
   46095 => x"ffffff",
   46096 => x"ffffff",
   46097 => x"ffffff",
   46098 => x"ffffff",
   46099 => x"ffffff",
   46100 => x"ffffff",
   46101 => x"ffffff",
   46102 => x"ffffff",
   46103 => x"ffffff",
   46104 => x"ffffff",
   46105 => x"ffffff",
   46106 => x"ffffff",
   46107 => x"ffffff",
   46108 => x"ffffff",
   46109 => x"ffffff",
   46110 => x"ffffff",
   46111 => x"ffffff",
   46112 => x"ffffff",
   46113 => x"ffffff",
   46114 => x"ffffff",
   46115 => x"ffffff",
   46116 => x"ffffff",
   46117 => x"ffffff",
   46118 => x"ffffff",
   46119 => x"ffffff",
   46120 => x"ffffff",
   46121 => x"ffffff",
   46122 => x"ffffff",
   46123 => x"ffffff",
   46124 => x"ffffff",
   46125 => x"ffffff",
   46126 => x"ffffff",
   46127 => x"ffffff",
   46128 => x"ffffff",
   46129 => x"ffffff",
   46130 => x"ffffff",
   46131 => x"ffffff",
   46132 => x"ffffff",
   46133 => x"ffffff",
   46134 => x"ffffff",
   46135 => x"ffffff",
   46136 => x"ffffff",
   46137 => x"ffffff",
   46138 => x"ffffff",
   46139 => x"ffffff",
   46140 => x"ffffff",
   46141 => x"ffffff",
   46142 => x"ffffff",
   46143 => x"ffffff",
   46144 => x"ffffff",
   46145 => x"ffffff",
   46146 => x"ffffff",
   46147 => x"ffffff",
   46148 => x"ffffff",
   46149 => x"fffa95",
   46150 => x"abffff",
   46151 => x"ffffff",
   46152 => x"ffffff",
   46153 => x"ffffff",
   46154 => x"ffffff",
   46155 => x"ffffff",
   46156 => x"ffffff",
   46157 => x"ffffff",
   46158 => x"ffffff",
   46159 => x"ffffff",
   46160 => x"ffffff",
   46161 => x"ffffff",
   46162 => x"ffffff",
   46163 => x"ffffff",
   46164 => x"ffffff",
   46165 => x"ffffff",
   46166 => x"ffffff",
   46167 => x"ffffff",
   46168 => x"ffffff",
   46169 => x"ffffff",
   46170 => x"ffffff",
   46171 => x"ffffff",
   46172 => x"ffffff",
   46173 => x"ffffff",
   46174 => x"ffffff",
   46175 => x"ffffff",
   46176 => x"ffffff",
   46177 => x"ffffff",
   46178 => x"ffffff",
   46179 => x"ffffff",
   46180 => x"ffffff",
   46181 => x"ffffff",
   46182 => x"ffffff",
   46183 => x"ffffff",
   46184 => x"ffffff",
   46185 => x"ffffff",
   46186 => x"ffffff",
   46187 => x"ffffff",
   46188 => x"ffffff",
   46189 => x"ffffff",
   46190 => x"ffffff",
   46191 => x"ffffff",
   46192 => x"ffffff",
   46193 => x"ffffff",
   46194 => x"ffffff",
   46195 => x"ffffff",
   46196 => x"ffffff",
   46197 => x"ffffff",
   46198 => x"ffffff",
   46199 => x"ffffff",
   46200 => x"ffffff",
   46201 => x"ffffff",
   46202 => x"ffffff",
   46203 => x"ffffff",
   46204 => x"ffffff",
   46205 => x"ffffff",
   46206 => x"ffffff",
   46207 => x"ffffff",
   46208 => x"ffffff",
   46209 => x"ffffff",
   46210 => x"ffffff",
   46211 => x"ffffff",
   46212 => x"ffffff",
   46213 => x"ffffff",
   46214 => x"ffffff",
   46215 => x"ffffff",
   46216 => x"ffffff",
   46217 => x"ffffff",
   46218 => x"ffffff",
   46219 => x"ffffff",
   46220 => x"ffffff",
   46221 => x"ffffff",
   46222 => x"ffffff",
   46223 => x"ffffff",
   46224 => x"ffffff",
   46225 => x"ffffff",
   46226 => x"ffffff",
   46227 => x"ffffff",
   46228 => x"ffffff",
   46229 => x"ffffff",
   46230 => x"ffffff",
   46231 => x"ffffff",
   46232 => x"ffffff",
   46233 => x"ffffff",
   46234 => x"ffffff",
   46235 => x"ffffff",
   46236 => x"ffffff",
   46237 => x"ffffff",
   46238 => x"ffffff",
   46239 => x"ffffff",
   46240 => x"ffffff",
   46241 => x"ffffff",
   46242 => x"ffffff",
   46243 => x"ffffff",
   46244 => x"ffffff",
   46245 => x"ffffff",
   46246 => x"ffffff",
   46247 => x"ffffff",
   46248 => x"ffffff",
   46249 => x"ffffff",
   46250 => x"ffffff",
   46251 => x"ffffff",
   46252 => x"ffffff",
   46253 => x"ffffff",
   46254 => x"ffffff",
   46255 => x"ffffff",
   46256 => x"ffffff",
   46257 => x"ffffff",
   46258 => x"ffffff",
   46259 => x"ffffff",
   46260 => x"ffffff",
   46261 => x"ffffff",
   46262 => x"ffffff",
   46263 => x"ffffff",
   46264 => x"ffffff",
   46265 => x"ffffff",
   46266 => x"ffffff",
   46267 => x"ffffff",
   46268 => x"ffffff",
   46269 => x"ffffff",
   46270 => x"ffffff",
   46271 => x"ffffff",
   46272 => x"ffffff",
   46273 => x"ffffff",
   46274 => x"ffffff",
   46275 => x"ffffff",
   46276 => x"ffffff",
   46277 => x"ffffff",
   46278 => x"ffffff",
   46279 => x"ffffff",
   46280 => x"ffffff",
   46281 => x"ffffff",
   46282 => x"ffffff",
   46283 => x"ffffff",
   46284 => x"ffffff",
   46285 => x"ffffff",
   46286 => x"ffffff",
   46287 => x"ffffff",
   46288 => x"ffffff",
   46289 => x"ffffff",
   46290 => x"ffffff",
   46291 => x"ffffff",
   46292 => x"ffffff",
   46293 => x"ffffff",
   46294 => x"ffffff",
   46295 => x"ffffff",
   46296 => x"ffffff",
   46297 => x"ffffff",
   46298 => x"ffffff",
   46299 => x"ffffff",
   46300 => x"ffffff",
   46301 => x"ffffff",
   46302 => x"ffffff",
   46303 => x"ffffff",
   46304 => x"ffffff",
   46305 => x"ffffff",
   46306 => x"ffffff",
   46307 => x"ffffff",
   46308 => x"ffffff",
   46309 => x"fffa95",
   46310 => x"abffff",
   46311 => x"ffffff",
   46312 => x"ffffff",
   46313 => x"ffffff",
   46314 => x"ffffff",
   46315 => x"ffffff",
   46316 => x"ffffff",
   46317 => x"ffffff",
   46318 => x"ffffff",
   46319 => x"ffffff",
   46320 => x"ffffff",
   46321 => x"ffffff",
   46322 => x"ffffff",
   46323 => x"ffffff",
   46324 => x"ffffff",
   46325 => x"ffffff",
   46326 => x"ffffff",
   46327 => x"ffffff",
   46328 => x"ffffff",
   46329 => x"ffffff",
   46330 => x"ffffff",
   46331 => x"ffffff",
   46332 => x"ffffff",
   46333 => x"ffffff",
   46334 => x"ffffff",
   46335 => x"ffffff",
   46336 => x"ffffff",
   46337 => x"ffffff",
   46338 => x"ffffff",
   46339 => x"ffffff",
   46340 => x"ffffff",
   46341 => x"ffffff",
   46342 => x"ffffff",
   46343 => x"ffffff",
   46344 => x"ffffff",
   46345 => x"ffffff",
   46346 => x"ffffff",
   46347 => x"ffffff",
   46348 => x"ffffff",
   46349 => x"ffffff",
   46350 => x"ffffff",
   46351 => x"ffffff",
   46352 => x"ffffff",
   46353 => x"ffffff",
   46354 => x"ffffff",
   46355 => x"ffffff",
   46356 => x"ffffff",
   46357 => x"ffffff",
   46358 => x"ffffff",
   46359 => x"ffffff",
   46360 => x"ffffff",
   46361 => x"ffffff",
   46362 => x"ffffff",
   46363 => x"ffffff",
   46364 => x"ffffff",
   46365 => x"ffffff",
   46366 => x"ffffff",
   46367 => x"ffffff",
   46368 => x"ffffff",
   46369 => x"ffffff",
   46370 => x"ffffff",
   46371 => x"ffffff",
   46372 => x"ffffff",
   46373 => x"ffffff",
   46374 => x"ffffff",
   46375 => x"ffffff",
   46376 => x"ffffff",
   46377 => x"ffffff",
   46378 => x"ffffff",
   46379 => x"ffffff",
   46380 => x"ffffff",
   46381 => x"ffffff",
   46382 => x"ffffff",
   46383 => x"ffffff",
   46384 => x"ffffff",
   46385 => x"ffffff",
   46386 => x"ffffff",
   46387 => x"ffffff",
   46388 => x"ffffff",
   46389 => x"ffffff",
   46390 => x"ffffff",
   46391 => x"ffffff",
   46392 => x"ffffff",
   46393 => x"ffffff",
   46394 => x"ffffff",
   46395 => x"ffffff",
   46396 => x"ffffff",
   46397 => x"ffffff",
   46398 => x"ffffff",
   46399 => x"ffffff",
   46400 => x"ffffff",
   46401 => x"ffffff",
   46402 => x"ffffff",
   46403 => x"ffffff",
   46404 => x"ffffff",
   46405 => x"ffffff",
   46406 => x"ffffff",
   46407 => x"ffffff",
   46408 => x"ffffff",
   46409 => x"ffffff",
   46410 => x"ffffff",
   46411 => x"ffffff",
   46412 => x"ffffff",
   46413 => x"ffffff",
   46414 => x"ffffff",
   46415 => x"ffffff",
   46416 => x"ffffff",
   46417 => x"ffffff",
   46418 => x"ffffff",
   46419 => x"ffffff",
   46420 => x"ffffff",
   46421 => x"ffffff",
   46422 => x"ffffff",
   46423 => x"ffffff",
   46424 => x"ffffff",
   46425 => x"ffffff",
   46426 => x"ffffff",
   46427 => x"ffffff",
   46428 => x"ffffff",
   46429 => x"ffffff",
   46430 => x"ffffff",
   46431 => x"ffffff",
   46432 => x"ffffff",
   46433 => x"ffffff",
   46434 => x"ffffff",
   46435 => x"ffffff",
   46436 => x"ffffff",
   46437 => x"ffffff",
   46438 => x"ffffff",
   46439 => x"ffffff",
   46440 => x"ffffff",
   46441 => x"ffffff",
   46442 => x"ffffff",
   46443 => x"ffffff",
   46444 => x"ffffff",
   46445 => x"ffffff",
   46446 => x"ffffff",
   46447 => x"ffffff",
   46448 => x"ffffff",
   46449 => x"ffffff",
   46450 => x"ffffff",
   46451 => x"ffffff",
   46452 => x"ffffff",
   46453 => x"ffffff",
   46454 => x"ffffff",
   46455 => x"ffffff",
   46456 => x"ffffff",
   46457 => x"ffffff",
   46458 => x"ffffff",
   46459 => x"ffffff",
   46460 => x"ffffff",
   46461 => x"ffffff",
   46462 => x"ffffff",
   46463 => x"ffffff",
   46464 => x"ffffff",
   46465 => x"ffffff",
   46466 => x"ffffff",
   46467 => x"ffffff",
   46468 => x"ffffff",
   46469 => x"fffa95",
   46470 => x"abffff",
   46471 => x"ffffff",
   46472 => x"ffffff",
   46473 => x"ffffff",
   46474 => x"ffffff",
   46475 => x"ffffff",
   46476 => x"ffffff",
   46477 => x"ffffff",
   46478 => x"ffffff",
   46479 => x"ffffff",
   46480 => x"ffffff",
   46481 => x"ffffff",
   46482 => x"ffffff",
   46483 => x"ffffff",
   46484 => x"ffffff",
   46485 => x"ffffff",
   46486 => x"ffffff",
   46487 => x"ffffff",
   46488 => x"ffffff",
   46489 => x"ffffff",
   46490 => x"ffffff",
   46491 => x"ffffff",
   46492 => x"ffffff",
   46493 => x"ffffff",
   46494 => x"ffffff",
   46495 => x"ffffff",
   46496 => x"ffffff",
   46497 => x"ffffff",
   46498 => x"ffffff",
   46499 => x"ffffff",
   46500 => x"ffffff",
   46501 => x"ffffff",
   46502 => x"ffffff",
   46503 => x"ffffff",
   46504 => x"ffffff",
   46505 => x"ffffff",
   46506 => x"ffffff",
   46507 => x"ffffff",
   46508 => x"ffffff",
   46509 => x"ffffff",
   46510 => x"ffffff",
   46511 => x"ffffff",
   46512 => x"ffffff",
   46513 => x"ffffff",
   46514 => x"ffffff",
   46515 => x"ffffff",
   46516 => x"ffffff",
   46517 => x"ffffff",
   46518 => x"ffffff",
   46519 => x"ffffff",
   46520 => x"ffffff",
   46521 => x"ffffff",
   46522 => x"ffffff",
   46523 => x"ffffff",
   46524 => x"ffffff",
   46525 => x"ffffff",
   46526 => x"ffffff",
   46527 => x"ffffff",
   46528 => x"ffffff",
   46529 => x"ffffff",
   46530 => x"ffffff",
   46531 => x"ffffff",
   46532 => x"ffffff",
   46533 => x"ffffff",
   46534 => x"ffffff",
   46535 => x"ffffff",
   46536 => x"ffffff",
   46537 => x"ffffff",
   46538 => x"ffffff",
   46539 => x"ffffff",
   46540 => x"ffffff",
   46541 => x"ffffff",
   46542 => x"ffffff",
   46543 => x"ffffff",
   46544 => x"ffffff",
   46545 => x"ffffff",
   46546 => x"ffffff",
   46547 => x"ffffff",
   46548 => x"ffffff",
   46549 => x"ffffff",
   46550 => x"ffffff",
   46551 => x"ffffff",
   46552 => x"ffffff",
   46553 => x"ffffff",
   46554 => x"ffffff",
   46555 => x"ffffff",
   46556 => x"ffffff",
   46557 => x"ffffff",
   46558 => x"ffffff",
   46559 => x"ffffff",
   46560 => x"ffffff",
   46561 => x"ffffff",
   46562 => x"ffffff",
   46563 => x"ffffff",
   46564 => x"ffffff",
   46565 => x"ffffff",
   46566 => x"ffffff",
   46567 => x"ffffff",
   46568 => x"ffffff",
   46569 => x"ffffff",
   46570 => x"ffffff",
   46571 => x"ffffff",
   46572 => x"ffffff",
   46573 => x"ffffff",
   46574 => x"ffffff",
   46575 => x"ffffff",
   46576 => x"ffffff",
   46577 => x"ffffff",
   46578 => x"ffffff",
   46579 => x"ffffff",
   46580 => x"ffffff",
   46581 => x"ffffff",
   46582 => x"ffffff",
   46583 => x"ffffff",
   46584 => x"ffffff",
   46585 => x"ffffff",
   46586 => x"ffffff",
   46587 => x"ffffff",
   46588 => x"ffffff",
   46589 => x"ffffff",
   46590 => x"ffffff",
   46591 => x"ffffff",
   46592 => x"ffffff",
   46593 => x"ffffff",
   46594 => x"ffffff",
   46595 => x"ffffff",
   46596 => x"ffffff",
   46597 => x"ffffff",
   46598 => x"ffffff",
   46599 => x"ffffff",
   46600 => x"ffffff",
   46601 => x"ffffff",
   46602 => x"ffffff",
   46603 => x"ffffff",
   46604 => x"ffffff",
   46605 => x"ffffff",
   46606 => x"ffffff",
   46607 => x"ffffff",
   46608 => x"ffffff",
   46609 => x"ffffff",
   46610 => x"ffffff",
   46611 => x"ffffff",
   46612 => x"ffffff",
   46613 => x"ffffff",
   46614 => x"ffffff",
   46615 => x"ffffff",
   46616 => x"ffffff",
   46617 => x"ffffff",
   46618 => x"ffffff",
   46619 => x"ffffff",
   46620 => x"ffffff",
   46621 => x"ffffff",
   46622 => x"ffffff",
   46623 => x"ffffff",
   46624 => x"ffffff",
   46625 => x"ffffff",
   46626 => x"ffffff",
   46627 => x"ffffff",
   46628 => x"ffffff",
   46629 => x"fffa95",
   46630 => x"abffff",
   46631 => x"ffffff",
   46632 => x"ffffff",
   46633 => x"ffffff",
   46634 => x"ffffff",
   46635 => x"ffffff",
   46636 => x"ffffff",
   46637 => x"ffffff",
   46638 => x"ffffff",
   46639 => x"ffffff",
   46640 => x"ffffff",
   46641 => x"ffffff",
   46642 => x"ffffff",
   46643 => x"ffffff",
   46644 => x"ffffff",
   46645 => x"ffffff",
   46646 => x"ffffff",
   46647 => x"ffffff",
   46648 => x"ffffff",
   46649 => x"ffffff",
   46650 => x"ffffff",
   46651 => x"ffffff",
   46652 => x"ffffff",
   46653 => x"ffffff",
   46654 => x"ffffff",
   46655 => x"ffffff",
   46656 => x"ffffff",
   46657 => x"ffffff",
   46658 => x"ffffff",
   46659 => x"ffffff",
   46660 => x"ffffff",
   46661 => x"ffffff",
   46662 => x"ffffff",
   46663 => x"ffffff",
   46664 => x"ffffff",
   46665 => x"ffffff",
   46666 => x"ffffff",
   46667 => x"ffffff",
   46668 => x"ffffff",
   46669 => x"ffffff",
   46670 => x"ffffff",
   46671 => x"ffffff",
   46672 => x"ffffff",
   46673 => x"ffffff",
   46674 => x"ffffff",
   46675 => x"ffffff",
   46676 => x"ffffff",
   46677 => x"ffffff",
   46678 => x"ffffff",
   46679 => x"ffffff",
   46680 => x"ffffff",
   46681 => x"ffffff",
   46682 => x"ffffff",
   46683 => x"ffffff",
   46684 => x"ffffff",
   46685 => x"ffffff",
   46686 => x"ffffff",
   46687 => x"ffffff",
   46688 => x"ffffff",
   46689 => x"ffffff",
   46690 => x"ffffff",
   46691 => x"ffffff",
   46692 => x"ffffff",
   46693 => x"ffffff",
   46694 => x"ffffff",
   46695 => x"ffffff",
   46696 => x"ffffff",
   46697 => x"ffffff",
   46698 => x"ffffff",
   46699 => x"ffffff",
   46700 => x"ffffff",
   46701 => x"ffffff",
   46702 => x"ffffff",
   46703 => x"ffffff",
   46704 => x"ffffff",
   46705 => x"ffffff",
   46706 => x"ffffff",
   46707 => x"ffffff",
   46708 => x"ffffff",
   46709 => x"ffffff",
   46710 => x"ffffff",
   46711 => x"ffffff",
   46712 => x"ffffff",
   46713 => x"ffffff",
   46714 => x"ffffff",
   46715 => x"ffffff",
   46716 => x"ffffff",
   46717 => x"ffffff",
   46718 => x"ffffff",
   46719 => x"ffffff",
   46720 => x"ffffff",
   46721 => x"ffffff",
   46722 => x"ffffff",
   46723 => x"ffffff",
   46724 => x"ffffff",
   46725 => x"ffffff",
   46726 => x"ffffff",
   46727 => x"ffffff",
   46728 => x"ffffff",
   46729 => x"ffffff",
   46730 => x"ffffff",
   46731 => x"ffffff",
   46732 => x"ffffff",
   46733 => x"ffffff",
   46734 => x"ffffff",
   46735 => x"ffffff",
   46736 => x"ffffff",
   46737 => x"ffffff",
   46738 => x"ffffff",
   46739 => x"ffffff",
   46740 => x"ffffff",
   46741 => x"ffffff",
   46742 => x"ffffff",
   46743 => x"ffffff",
   46744 => x"ffffff",
   46745 => x"ffffff",
   46746 => x"ffffff",
   46747 => x"ffffff",
   46748 => x"ffffff",
   46749 => x"ffffff",
   46750 => x"ffffff",
   46751 => x"ffffff",
   46752 => x"ffffff",
   46753 => x"ffffff",
   46754 => x"ffffff",
   46755 => x"ffffff",
   46756 => x"ffffff",
   46757 => x"ffffff",
   46758 => x"ffffff",
   46759 => x"ffffff",
   46760 => x"ffffff",
   46761 => x"ffffff",
   46762 => x"ffffff",
   46763 => x"ffffff",
   46764 => x"ffffff",
   46765 => x"ffffff",
   46766 => x"ffffff",
   46767 => x"ffffff",
   46768 => x"ffffff",
   46769 => x"ffffff",
   46770 => x"ffffff",
   46771 => x"ffffff",
   46772 => x"ffffff",
   46773 => x"ffffff",
   46774 => x"ffffff",
   46775 => x"ffffff",
   46776 => x"ffffff",
   46777 => x"ffffff",
   46778 => x"ffffff",
   46779 => x"ffffff",
   46780 => x"ffffff",
   46781 => x"ffffff",
   46782 => x"ffffff",
   46783 => x"ffffff",
   46784 => x"ffffff",
   46785 => x"ffffff",
   46786 => x"ffffff",
   46787 => x"ffffff",
   46788 => x"ffffff",
   46789 => x"fffa95",
   46790 => x"abffff",
   46791 => x"ffffff",
   46792 => x"ffffff",
   46793 => x"ffffff",
   46794 => x"ffffff",
   46795 => x"ffffff",
   46796 => x"ffffff",
   46797 => x"ffffff",
   46798 => x"ffffff",
   46799 => x"ffffff",
   46800 => x"ffffff",
   46801 => x"ffffff",
   46802 => x"ffffff",
   46803 => x"ffffff",
   46804 => x"ffffff",
   46805 => x"ffffff",
   46806 => x"ffffff",
   46807 => x"ffffff",
   46808 => x"ffffff",
   46809 => x"ffffff",
   46810 => x"ffffff",
   46811 => x"ffffff",
   46812 => x"ffffff",
   46813 => x"ffffff",
   46814 => x"ffffff",
   46815 => x"ffffff",
   46816 => x"ffffff",
   46817 => x"ffffff",
   46818 => x"ffffff",
   46819 => x"ffffff",
   46820 => x"ffffff",
   46821 => x"ffffff",
   46822 => x"ffffff",
   46823 => x"ffffff",
   46824 => x"ffffff",
   46825 => x"ffffff",
   46826 => x"ffffff",
   46827 => x"ffffff",
   46828 => x"ffffff",
   46829 => x"ffffff",
   46830 => x"ffffff",
   46831 => x"ffffff",
   46832 => x"ffffff",
   46833 => x"ffffff",
   46834 => x"ffffff",
   46835 => x"ffffff",
   46836 => x"ffffff",
   46837 => x"ffffff",
   46838 => x"ffffff",
   46839 => x"ffffff",
   46840 => x"ffffff",
   46841 => x"ffffff",
   46842 => x"ffffff",
   46843 => x"ffffff",
   46844 => x"ffffff",
   46845 => x"ffffff",
   46846 => x"ffffff",
   46847 => x"ffffff",
   46848 => x"ffffff",
   46849 => x"ffffff",
   46850 => x"ffffff",
   46851 => x"ffffff",
   46852 => x"ffffff",
   46853 => x"ffffff",
   46854 => x"ffffff",
   46855 => x"ffffff",
   46856 => x"ffffff",
   46857 => x"ffffff",
   46858 => x"ffffff",
   46859 => x"ffffff",
   46860 => x"ffffff",
   46861 => x"ffffff",
   46862 => x"ffffff",
   46863 => x"ffffff",
   46864 => x"ffffff",
   46865 => x"ffffff",
   46866 => x"ffffff",
   46867 => x"ffffff",
   46868 => x"ffffff",
   46869 => x"ffffff",
   46870 => x"ffffff",
   46871 => x"ffffff",
   46872 => x"ffffff",
   46873 => x"ffffff",
   46874 => x"ffffff",
   46875 => x"ffffff",
   46876 => x"ffffff",
   46877 => x"ffffff",
   46878 => x"ffffff",
   46879 => x"ffffff",
   46880 => x"ffffff",
   46881 => x"ffffff",
   46882 => x"ffffff",
   46883 => x"ffffff",
   46884 => x"ffffff",
   46885 => x"ffffff",
   46886 => x"ffffff",
   46887 => x"ffffff",
   46888 => x"ffffff",
   46889 => x"ffffff",
   46890 => x"ffffff",
   46891 => x"ffffff",
   46892 => x"ffffff",
   46893 => x"ffffff",
   46894 => x"ffffff",
   46895 => x"ffffff",
   46896 => x"ffffff",
   46897 => x"ffffff",
   46898 => x"ffffff",
   46899 => x"ffffff",
   46900 => x"ffffff",
   46901 => x"ffffff",
   46902 => x"ffffff",
   46903 => x"ffffff",
   46904 => x"ffffff",
   46905 => x"ffffff",
   46906 => x"ffffff",
   46907 => x"ffffff",
   46908 => x"ffffff",
   46909 => x"ffffff",
   46910 => x"ffffff",
   46911 => x"ffffff",
   46912 => x"ffffff",
   46913 => x"ffffff",
   46914 => x"ffffff",
   46915 => x"ffffff",
   46916 => x"ffffff",
   46917 => x"ffffff",
   46918 => x"ffffff",
   46919 => x"ffffff",
   46920 => x"ffffff",
   46921 => x"ffffff",
   46922 => x"ffffff",
   46923 => x"ffffff",
   46924 => x"ffffff",
   46925 => x"ffffff",
   46926 => x"ffffff",
   46927 => x"ffffff",
   46928 => x"ffffff",
   46929 => x"ffffff",
   46930 => x"ffffff",
   46931 => x"ffffff",
   46932 => x"ffffff",
   46933 => x"ffffff",
   46934 => x"ffffff",
   46935 => x"ffffff",
   46936 => x"ffffff",
   46937 => x"ffffff",
   46938 => x"ffffff",
   46939 => x"ffffff",
   46940 => x"ffffff",
   46941 => x"ffffff",
   46942 => x"ffffff",
   46943 => x"ffffff",
   46944 => x"ffffff",
   46945 => x"ffffff",
   46946 => x"ffffff",
   46947 => x"ffffff",
   46948 => x"ffffff",
   46949 => x"fffa95",
   46950 => x"abffff",
   46951 => x"ffffff",
   46952 => x"ffffff",
   46953 => x"ffffff",
   46954 => x"ffffff",
   46955 => x"ffffff",
   46956 => x"ffffff",
   46957 => x"ffffff",
   46958 => x"ffffff",
   46959 => x"ffffff",
   46960 => x"ffffff",
   46961 => x"ffffff",
   46962 => x"ffffff",
   46963 => x"ffffff",
   46964 => x"ffffff",
   46965 => x"ffffff",
   46966 => x"ffffff",
   46967 => x"ffffff",
   46968 => x"ffffff",
   46969 => x"ffffff",
   46970 => x"ffffff",
   46971 => x"ffffff",
   46972 => x"ffffff",
   46973 => x"ffffff",
   46974 => x"ffffff",
   46975 => x"ffffff",
   46976 => x"ffffff",
   46977 => x"ffffff",
   46978 => x"ffffff",
   46979 => x"ffffff",
   46980 => x"ffffff",
   46981 => x"ffffff",
   46982 => x"ffffff",
   46983 => x"ffffff",
   46984 => x"ffffff",
   46985 => x"ffffff",
   46986 => x"ffffff",
   46987 => x"ffffff",
   46988 => x"ffffff",
   46989 => x"ffffff",
   46990 => x"ffffff",
   46991 => x"ffffff",
   46992 => x"ffffff",
   46993 => x"ffffff",
   46994 => x"ffffff",
   46995 => x"ffffff",
   46996 => x"ffffff",
   46997 => x"ffffff",
   46998 => x"ffffff",
   46999 => x"ffffff",
   47000 => x"ffffff",
   47001 => x"ffffff",
   47002 => x"ffffff",
   47003 => x"ffffff",
   47004 => x"ffffff",
   47005 => x"ffffff",
   47006 => x"ffffff",
   47007 => x"ffffff",
   47008 => x"ffffff",
   47009 => x"ffffff",
   47010 => x"ffffff",
   47011 => x"ffffff",
   47012 => x"ffffff",
   47013 => x"ffffff",
   47014 => x"ffffff",
   47015 => x"ffffff",
   47016 => x"ffffff",
   47017 => x"ffffff",
   47018 => x"ffffff",
   47019 => x"ffffff",
   47020 => x"ffffff",
   47021 => x"ffffff",
   47022 => x"ffffff",
   47023 => x"ffffff",
   47024 => x"ffffff",
   47025 => x"ffffff",
   47026 => x"ffffff",
   47027 => x"ffffff",
   47028 => x"ffffff",
   47029 => x"ffffff",
   47030 => x"ffffff",
   47031 => x"ffffff",
   47032 => x"ffffff",
   47033 => x"ffffff",
   47034 => x"ffffff",
   47035 => x"ffffff",
   47036 => x"ffffff",
   47037 => x"ffffff",
   47038 => x"ffffff",
   47039 => x"ffffff",
   47040 => x"ffffff",
   47041 => x"ffffff",
   47042 => x"ffffff",
   47043 => x"ffffff",
   47044 => x"ffffff",
   47045 => x"ffffff",
   47046 => x"ffffff",
   47047 => x"ffffff",
   47048 => x"ffffff",
   47049 => x"ffffff",
   47050 => x"ffffff",
   47051 => x"ffffff",
   47052 => x"ffffff",
   47053 => x"ffffff",
   47054 => x"ffffff",
   47055 => x"ffffff",
   47056 => x"ffffff",
   47057 => x"ffffff",
   47058 => x"ffffff",
   47059 => x"ffffff",
   47060 => x"ffffff",
   47061 => x"ffffff",
   47062 => x"ffffff",
   47063 => x"ffffff",
   47064 => x"ffffff",
   47065 => x"ffffff",
   47066 => x"ffffff",
   47067 => x"ffffff",
   47068 => x"ffffff",
   47069 => x"ffffff",
   47070 => x"ffffff",
   47071 => x"ffffff",
   47072 => x"ffffff",
   47073 => x"ffffff",
   47074 => x"ffffff",
   47075 => x"ffffff",
   47076 => x"ffffff",
   47077 => x"ffffff",
   47078 => x"ffffff",
   47079 => x"ffffff",
   47080 => x"ffffff",
   47081 => x"ffffff",
   47082 => x"ffffff",
   47083 => x"ffffff",
   47084 => x"ffffff",
   47085 => x"ffffff",
   47086 => x"ffffff",
   47087 => x"ffffff",
   47088 => x"ffffff",
   47089 => x"ffffff",
   47090 => x"ffffff",
   47091 => x"ffffff",
   47092 => x"ffffff",
   47093 => x"ffffff",
   47094 => x"ffffff",
   47095 => x"ffffff",
   47096 => x"ffffff",
   47097 => x"ffffff",
   47098 => x"ffffff",
   47099 => x"ffffff",
   47100 => x"ffffff",
   47101 => x"ffffff",
   47102 => x"ffffff",
   47103 => x"ffffff",
   47104 => x"ffffff",
   47105 => x"ffffff",
   47106 => x"ffffff",
   47107 => x"ffffff",
   47108 => x"ffffff",
   47109 => x"fffa95",
   47110 => x"abffff",
   47111 => x"ffffff",
   47112 => x"ffffff",
   47113 => x"ffffff",
   47114 => x"ffffff",
   47115 => x"ffffff",
   47116 => x"ffffff",
   47117 => x"ffffff",
   47118 => x"ffffff",
   47119 => x"ffffff",
   47120 => x"ffffff",
   47121 => x"ffffff",
   47122 => x"ffffff",
   47123 => x"ffffff",
   47124 => x"ffffff",
   47125 => x"ffffff",
   47126 => x"ffffff",
   47127 => x"ffffff",
   47128 => x"ffffff",
   47129 => x"ffffff",
   47130 => x"ffffff",
   47131 => x"ffffff",
   47132 => x"ffffff",
   47133 => x"ffffff",
   47134 => x"ffffff",
   47135 => x"ffffff",
   47136 => x"ffffff",
   47137 => x"ffffff",
   47138 => x"ffffff",
   47139 => x"ffffff",
   47140 => x"ffffff",
   47141 => x"ffffff",
   47142 => x"ffffff",
   47143 => x"ffffff",
   47144 => x"ffffff",
   47145 => x"ffffff",
   47146 => x"ffffff",
   47147 => x"ffffff",
   47148 => x"ffffff",
   47149 => x"ffffff",
   47150 => x"ffffff",
   47151 => x"ffffff",
   47152 => x"ffffff",
   47153 => x"ffffff",
   47154 => x"ffffff",
   47155 => x"ffffff",
   47156 => x"ffffff",
   47157 => x"ffffff",
   47158 => x"ffffff",
   47159 => x"ffffff",
   47160 => x"ffffff",
   47161 => x"ffffff",
   47162 => x"ffffff",
   47163 => x"ffffff",
   47164 => x"ffffff",
   47165 => x"ffffff",
   47166 => x"ffffff",
   47167 => x"ffffff",
   47168 => x"ffffff",
   47169 => x"ffffff",
   47170 => x"ffffff",
   47171 => x"ffffff",
   47172 => x"ffffff",
   47173 => x"ffffff",
   47174 => x"ffffff",
   47175 => x"ffffff",
   47176 => x"ffffff",
   47177 => x"ffffff",
   47178 => x"ffffff",
   47179 => x"ffffff",
   47180 => x"ffffff",
   47181 => x"ffffff",
   47182 => x"ffffff",
   47183 => x"ffffff",
   47184 => x"ffffff",
   47185 => x"ffffff",
   47186 => x"ffffff",
   47187 => x"ffffff",
   47188 => x"ffffff",
   47189 => x"ffffff",
   47190 => x"ffffff",
   47191 => x"ffffff",
   47192 => x"ffffff",
   47193 => x"ffffff",
   47194 => x"ffffff",
   47195 => x"ffffff",
   47196 => x"ffffff",
   47197 => x"ffffff",
   47198 => x"ffffff",
   47199 => x"ffffff",
   47200 => x"ffffff",
   47201 => x"ffffff",
   47202 => x"ffffff",
   47203 => x"ffffff",
   47204 => x"ffffff",
   47205 => x"ffffff",
   47206 => x"ffffff",
   47207 => x"ffffff",
   47208 => x"ffffff",
   47209 => x"ffffff",
   47210 => x"ffffff",
   47211 => x"ffffff",
   47212 => x"ffffff",
   47213 => x"ffffff",
   47214 => x"ffffff",
   47215 => x"ffffff",
   47216 => x"ffffff",
   47217 => x"ffffff",
   47218 => x"ffffff",
   47219 => x"ffffff",
   47220 => x"ffffff",
   47221 => x"ffffff",
   47222 => x"ffffff",
   47223 => x"ffffff",
   47224 => x"ffffff",
   47225 => x"ffffff",
   47226 => x"ffffff",
   47227 => x"ffffff",
   47228 => x"ffffff",
   47229 => x"ffffff",
   47230 => x"ffffff",
   47231 => x"ffffff",
   47232 => x"ffffff",
   47233 => x"ffffff",
   47234 => x"ffffff",
   47235 => x"ffffff",
   47236 => x"ffffff",
   47237 => x"ffffff",
   47238 => x"ffffff",
   47239 => x"ffffff",
   47240 => x"ffffff",
   47241 => x"ffffff",
   47242 => x"ffffff",
   47243 => x"ffffff",
   47244 => x"ffffff",
   47245 => x"ffffff",
   47246 => x"ffffff",
   47247 => x"ffffff",
   47248 => x"ffffff",
   47249 => x"ffffff",
   47250 => x"ffffff",
   47251 => x"ffffff",
   47252 => x"ffffff",
   47253 => x"ffffff",
   47254 => x"ffffff",
   47255 => x"ffffff",
   47256 => x"ffffff",
   47257 => x"ffffff",
   47258 => x"ffffff",
   47259 => x"ffffff",
   47260 => x"ffffff",
   47261 => x"ffffff",
   47262 => x"ffffff",
   47263 => x"ffffff",
   47264 => x"ffffff",
   47265 => x"ffffff",
   47266 => x"ffffff",
   47267 => x"ffffff",
   47268 => x"ffffff",
   47269 => x"fffa95",
   47270 => x"abffff",
   47271 => x"ffffff",
   47272 => x"ffffff",
   47273 => x"ffffff",
   47274 => x"ffffff",
   47275 => x"ffffff",
   47276 => x"ffffff",
   47277 => x"ffffff",
   47278 => x"ffffff",
   47279 => x"ffffff",
   47280 => x"ffffff",
   47281 => x"ffffff",
   47282 => x"ffffff",
   47283 => x"ffffff",
   47284 => x"ffffff",
   47285 => x"ffffff",
   47286 => x"ffffff",
   47287 => x"ffffff",
   47288 => x"ffffff",
   47289 => x"ffffff",
   47290 => x"ffffff",
   47291 => x"ffffff",
   47292 => x"ffffff",
   47293 => x"ffffff",
   47294 => x"ffffff",
   47295 => x"ffffff",
   47296 => x"ffffff",
   47297 => x"ffffff",
   47298 => x"ffffff",
   47299 => x"ffffff",
   47300 => x"ffffff",
   47301 => x"ffffff",
   47302 => x"ffffff",
   47303 => x"ffffff",
   47304 => x"ffffff",
   47305 => x"ffffff",
   47306 => x"ffffff",
   47307 => x"ffffff",
   47308 => x"ffffff",
   47309 => x"ffffff",
   47310 => x"ffffff",
   47311 => x"ffffff",
   47312 => x"ffffff",
   47313 => x"ffffff",
   47314 => x"ffffff",
   47315 => x"ffffff",
   47316 => x"ffffff",
   47317 => x"ffffff",
   47318 => x"ffffff",
   47319 => x"ffffff",
   47320 => x"ffffff",
   47321 => x"ffffff",
   47322 => x"ffffff",
   47323 => x"ffffff",
   47324 => x"ffffff",
   47325 => x"ffffff",
   47326 => x"ffffff",
   47327 => x"ffffff",
   47328 => x"ffffff",
   47329 => x"ffffff",
   47330 => x"ffffff",
   47331 => x"ffffff",
   47332 => x"ffffff",
   47333 => x"ffffff",
   47334 => x"ffffff",
   47335 => x"ffffff",
   47336 => x"ffffff",
   47337 => x"ffffff",
   47338 => x"ffffff",
   47339 => x"ffffff",
   47340 => x"ffffff",
   47341 => x"ffffff",
   47342 => x"ffffff",
   47343 => x"ffffff",
   47344 => x"ffffff",
   47345 => x"ffffff",
   47346 => x"ffffff",
   47347 => x"ffffff",
   47348 => x"ffffff",
   47349 => x"ffffff",
   47350 => x"ffffff",
   47351 => x"ffffff",
   47352 => x"ffffff",
   47353 => x"ffffff",
   47354 => x"ffffff",
   47355 => x"ffffff",
   47356 => x"ffffff",
   47357 => x"ffffff",
   47358 => x"ffffff",
   47359 => x"ffffff",
   47360 => x"ffffff",
   47361 => x"ffffff",
   47362 => x"ffffff",
   47363 => x"ffffff",
   47364 => x"ffffff",
   47365 => x"ffffff",
   47366 => x"ffffff",
   47367 => x"ffffff",
   47368 => x"ffffff",
   47369 => x"ffffff",
   47370 => x"ffffff",
   47371 => x"ffffff",
   47372 => x"ffffff",
   47373 => x"ffffff",
   47374 => x"ffffff",
   47375 => x"ffffff",
   47376 => x"ffffff",
   47377 => x"ffffff",
   47378 => x"ffffff",
   47379 => x"ffffff",
   47380 => x"ffffff",
   47381 => x"ffffff",
   47382 => x"ffffff",
   47383 => x"ffffff",
   47384 => x"ffffff",
   47385 => x"ffffff",
   47386 => x"ffffff",
   47387 => x"ffffff",
   47388 => x"ffffff",
   47389 => x"ffffff",
   47390 => x"ffffff",
   47391 => x"ffffff",
   47392 => x"ffffff",
   47393 => x"ffffff",
   47394 => x"ffffff",
   47395 => x"ffffff",
   47396 => x"ffffff",
   47397 => x"ffffff",
   47398 => x"ffffff",
   47399 => x"ffffff",
   47400 => x"ffffff",
   47401 => x"ffffff",
   47402 => x"ffffff",
   47403 => x"ffffff",
   47404 => x"ffffff",
   47405 => x"ffffff",
   47406 => x"ffffff",
   47407 => x"ffffff",
   47408 => x"ffffff",
   47409 => x"ffffff",
   47410 => x"ffffff",
   47411 => x"ffffff",
   47412 => x"ffffff",
   47413 => x"ffffff",
   47414 => x"ffffff",
   47415 => x"ffffff",
   47416 => x"ffffff",
   47417 => x"ffffff",
   47418 => x"ffffff",
   47419 => x"ffffff",
   47420 => x"ffffff",
   47421 => x"ffffff",
   47422 => x"ffffff",
   47423 => x"ffffff",
   47424 => x"ffffff",
   47425 => x"ffffff",
   47426 => x"ffffff",
   47427 => x"ffffff",
   47428 => x"ffffff",
   47429 => x"fffa95",
   47430 => x"abffff",
   47431 => x"ffffff",
   47432 => x"ffffff",
   47433 => x"ffffff",
   47434 => x"ffffff",
   47435 => x"ffffff",
   47436 => x"ffffff",
   47437 => x"ffffff",
   47438 => x"ffffff",
   47439 => x"ffffff",
   47440 => x"ffffff",
   47441 => x"ffffff",
   47442 => x"ffffff",
   47443 => x"ffffff",
   47444 => x"ffffff",
   47445 => x"ffffff",
   47446 => x"ffffff",
   47447 => x"ffffff",
   47448 => x"ffffff",
   47449 => x"ffffff",
   47450 => x"ffffff",
   47451 => x"ffffff",
   47452 => x"ffffff",
   47453 => x"ffffff",
   47454 => x"ffffff",
   47455 => x"ffffff",
   47456 => x"ffffff",
   47457 => x"ffffff",
   47458 => x"ffffff",
   47459 => x"ffffff",
   47460 => x"ffffff",
   47461 => x"ffffff",
   47462 => x"ffffff",
   47463 => x"ffffff",
   47464 => x"ffffff",
   47465 => x"ffffff",
   47466 => x"ffffff",
   47467 => x"ffffff",
   47468 => x"ffffff",
   47469 => x"ffffff",
   47470 => x"ffffff",
   47471 => x"ffffff",
   47472 => x"ffffff",
   47473 => x"ffffff",
   47474 => x"ffffff",
   47475 => x"ffffff",
   47476 => x"ffffff",
   47477 => x"ffffff",
   47478 => x"ffffff",
   47479 => x"ffffff",
   47480 => x"ffffff",
   47481 => x"ffffff",
   47482 => x"ffffff",
   47483 => x"ffffff",
   47484 => x"ffffff",
   47485 => x"ffffff",
   47486 => x"ffffff",
   47487 => x"ffffff",
   47488 => x"ffffff",
   47489 => x"ffffff",
   47490 => x"ffffff",
   47491 => x"ffffff",
   47492 => x"ffffff",
   47493 => x"ffffff",
   47494 => x"ffffff",
   47495 => x"ffffff",
   47496 => x"ffffff",
   47497 => x"ffffff",
   47498 => x"ffffff",
   47499 => x"ffffff",
   47500 => x"ffffff",
   47501 => x"ffffff",
   47502 => x"ffffff",
   47503 => x"ffffff",
   47504 => x"ffffff",
   47505 => x"ffffff",
   47506 => x"ffffff",
   47507 => x"ffffff",
   47508 => x"ffffff",
   47509 => x"ffffff",
   47510 => x"ffffff",
   47511 => x"ffffff",
   47512 => x"ffffff",
   47513 => x"ffffff",
   47514 => x"ffffff",
   47515 => x"ffffff",
   47516 => x"ffffff",
   47517 => x"ffffff",
   47518 => x"ffffff",
   47519 => x"ffffff",
   47520 => x"ffffff",
   47521 => x"ffffff",
   47522 => x"ffffff",
   47523 => x"ffffff",
   47524 => x"ffffff",
   47525 => x"ffffff",
   47526 => x"ffffff",
   47527 => x"ffffff",
   47528 => x"ffffff",
   47529 => x"ffffff",
   47530 => x"ffffff",
   47531 => x"ffffff",
   47532 => x"ffffff",
   47533 => x"ffffff",
   47534 => x"ffffff",
   47535 => x"ffffff",
   47536 => x"ffffff",
   47537 => x"ffffff",
   47538 => x"ffffff",
   47539 => x"ffffff",
   47540 => x"ffffff",
   47541 => x"ffffff",
   47542 => x"ffffff",
   47543 => x"ffffff",
   47544 => x"ffffff",
   47545 => x"ffffff",
   47546 => x"ffffff",
   47547 => x"ffffff",
   47548 => x"ffffff",
   47549 => x"ffffff",
   47550 => x"ffffff",
   47551 => x"ffffff",
   47552 => x"ffffff",
   47553 => x"ffffff",
   47554 => x"ffffff",
   47555 => x"ffffff",
   47556 => x"ffffff",
   47557 => x"ffffff",
   47558 => x"ffffff",
   47559 => x"ffffff",
   47560 => x"ffffff",
   47561 => x"ffffff",
   47562 => x"ffffff",
   47563 => x"ffffff",
   47564 => x"ffffff",
   47565 => x"ffffff",
   47566 => x"ffffff",
   47567 => x"ffffff",
   47568 => x"ffffff",
   47569 => x"ffffff",
   47570 => x"ffffff",
   47571 => x"ffffff",
   47572 => x"ffffff",
   47573 => x"ffffff",
   47574 => x"ffffff",
   47575 => x"ffffff",
   47576 => x"ffffff",
   47577 => x"ffffff",
   47578 => x"ffffff",
   47579 => x"ffffff",
   47580 => x"ffffff",
   47581 => x"ffffff",
   47582 => x"ffffff",
   47583 => x"ffffff",
   47584 => x"ffffff",
   47585 => x"ffffff",
   47586 => x"ffffff",
   47587 => x"ffffff",
   47588 => x"ffffff",
   47589 => x"fffa95",
   47590 => x"abffff",
   47591 => x"ffffff",
   47592 => x"ffffff",
   47593 => x"ffffff",
   47594 => x"ffffff",
   47595 => x"ffffff",
   47596 => x"ffffff",
   47597 => x"ffffff",
   47598 => x"ffffff",
   47599 => x"ffffff",
   47600 => x"ffffff",
   47601 => x"ffffff",
   47602 => x"ffffff",
   47603 => x"ffffff",
   47604 => x"ffffff",
   47605 => x"ffffff",
   47606 => x"ffffff",
   47607 => x"ffffff",
   47608 => x"ffffff",
   47609 => x"ffffff",
   47610 => x"ffffff",
   47611 => x"ffffff",
   47612 => x"ffffff",
   47613 => x"ffffff",
   47614 => x"ffffff",
   47615 => x"ffffff",
   47616 => x"ffffff",
   47617 => x"ffffff",
   47618 => x"ffffff",
   47619 => x"ffffff",
   47620 => x"ffffff",
   47621 => x"ffffff",
   47622 => x"ffffff",
   47623 => x"ffffff",
   47624 => x"ffffff",
   47625 => x"ffffff",
   47626 => x"ffffff",
   47627 => x"ffffff",
   47628 => x"ffffff",
   47629 => x"ffffff",
   47630 => x"ffffff",
   47631 => x"ffffff",
   47632 => x"ffffff",
   47633 => x"ffffff",
   47634 => x"ffffff",
   47635 => x"ffffff",
   47636 => x"ffffff",
   47637 => x"ffffff",
   47638 => x"ffffff",
   47639 => x"ffffff",
   47640 => x"ffffff",
   47641 => x"ffffff",
   47642 => x"ffffff",
   47643 => x"ffffff",
   47644 => x"ffffff",
   47645 => x"ffffff",
   47646 => x"ffffff",
   47647 => x"ffffff",
   47648 => x"ffffff",
   47649 => x"ffffff",
   47650 => x"ffffff",
   47651 => x"ffffff",
   47652 => x"ffffff",
   47653 => x"ffffff",
   47654 => x"ffffff",
   47655 => x"ffffff",
   47656 => x"ffffff",
   47657 => x"ffffff",
   47658 => x"ffffff",
   47659 => x"ffffff",
   47660 => x"ffffff",
   47661 => x"ffffff",
   47662 => x"ffffff",
   47663 => x"ffffff",
   47664 => x"ffffff",
   47665 => x"ffffff",
   47666 => x"ffffff",
   47667 => x"ffffff",
   47668 => x"ffffff",
   47669 => x"ffffff",
   47670 => x"ffffff",
   47671 => x"ffffff",
   47672 => x"ffffff",
   47673 => x"ffffff",
   47674 => x"ffffff",
   47675 => x"ffffff",
   47676 => x"ffffff",
   47677 => x"ffffff",
   47678 => x"ffffff",
   47679 => x"ffffff",
   47680 => x"ffffff",
   47681 => x"ffffff",
   47682 => x"ffffff",
   47683 => x"ffffff",
   47684 => x"ffffff",
   47685 => x"ffffff",
   47686 => x"ffffff",
   47687 => x"ffffff",
   47688 => x"ffffff",
   47689 => x"ffffff",
   47690 => x"ffffff",
   47691 => x"ffffff",
   47692 => x"ffffff",
   47693 => x"ffffff",
   47694 => x"ffffff",
   47695 => x"ffffff",
   47696 => x"ffffff",
   47697 => x"ffffff",
   47698 => x"ffffff",
   47699 => x"ffffff",
   47700 => x"ffffff",
   47701 => x"ffffff",
   47702 => x"ffffff",
   47703 => x"ffffff",
   47704 => x"ffffff",
   47705 => x"ffffff",
   47706 => x"ffffff",
   47707 => x"ffffff",
   47708 => x"ffffff",
   47709 => x"ffffff",
   47710 => x"ffffff",
   47711 => x"ffffff",
   47712 => x"ffffff",
   47713 => x"ffffff",
   47714 => x"ffffff",
   47715 => x"ffffff",
   47716 => x"ffffff",
   47717 => x"ffffff",
   47718 => x"ffffff",
   47719 => x"ffffff",
   47720 => x"ffffff",
   47721 => x"ffffff",
   47722 => x"ffffff",
   47723 => x"ffffff",
   47724 => x"ffffff",
   47725 => x"ffffff",
   47726 => x"ffffff",
   47727 => x"ffffff",
   47728 => x"ffffff",
   47729 => x"ffffff",
   47730 => x"ffffff",
   47731 => x"ffffff",
   47732 => x"ffffff",
   47733 => x"ffffff",
   47734 => x"ffffff",
   47735 => x"ffffff",
   47736 => x"ffffff",
   47737 => x"ffffff",
   47738 => x"ffffff",
   47739 => x"ffffff",
   47740 => x"ffffff",
   47741 => x"ffffff",
   47742 => x"ffffff",
   47743 => x"ffffff",
   47744 => x"ffffff",
   47745 => x"ffffff",
   47746 => x"ffffff",
   47747 => x"ffffff",
   47748 => x"ffffff",
   47749 => x"fffa95",
   47750 => x"abffff",
   47751 => x"ffffff",
   47752 => x"ffffff",
   47753 => x"ffffff",
   47754 => x"ffffff",
   47755 => x"ffffff",
   47756 => x"ffffff",
   47757 => x"ffffff",
   47758 => x"ffffff",
   47759 => x"ffffff",
   47760 => x"ffffff",
   47761 => x"ffffff",
   47762 => x"ffffff",
   47763 => x"ffffff",
   47764 => x"ffffff",
   47765 => x"ffffff",
   47766 => x"ffffff",
   47767 => x"ffffff",
   47768 => x"ffffff",
   47769 => x"ffffff",
   47770 => x"ffffff",
   47771 => x"ffffff",
   47772 => x"ffffff",
   47773 => x"ffffff",
   47774 => x"ffffff",
   47775 => x"ffffff",
   47776 => x"ffffff",
   47777 => x"ffffff",
   47778 => x"ffffff",
   47779 => x"ffffff",
   47780 => x"ffffff",
   47781 => x"ffffff",
   47782 => x"ffffff",
   47783 => x"ffffff",
   47784 => x"ffffff",
   47785 => x"ffffff",
   47786 => x"ffffff",
   47787 => x"ffffff",
   47788 => x"ffffff",
   47789 => x"ffffff",
   47790 => x"ffffff",
   47791 => x"ffffff",
   47792 => x"ffffff",
   47793 => x"ffffff",
   47794 => x"ffffff",
   47795 => x"ffffff",
   47796 => x"ffffff",
   47797 => x"ffffff",
   47798 => x"ffffff",
   47799 => x"ffffff",
   47800 => x"ffffff",
   47801 => x"ffffff",
   47802 => x"ffffff",
   47803 => x"ffffff",
   47804 => x"ffffff",
   47805 => x"ffffff",
   47806 => x"ffffff",
   47807 => x"ffffff",
   47808 => x"ffffff",
   47809 => x"ffffff",
   47810 => x"ffffff",
   47811 => x"ffffff",
   47812 => x"ffffff",
   47813 => x"ffffff",
   47814 => x"ffffff",
   47815 => x"ffffff",
   47816 => x"ffffff",
   47817 => x"ffffff",
   47818 => x"ffffff",
   47819 => x"ffffff",
   47820 => x"ffffff",
   47821 => x"ffffff",
   47822 => x"ffffff",
   47823 => x"ffffff",
   47824 => x"ffffff",
   47825 => x"ffffff",
   47826 => x"ffffff",
   47827 => x"ffffff",
   47828 => x"ffffff",
   47829 => x"ffffff",
   47830 => x"ffffff",
   47831 => x"ffffff",
   47832 => x"ffffff",
   47833 => x"ffffff",
   47834 => x"ffffff",
   47835 => x"ffffff",
   47836 => x"ffffff",
   47837 => x"ffffff",
   47838 => x"ffffff",
   47839 => x"ffffff",
   47840 => x"ffffff",
   47841 => x"ffffff",
   47842 => x"ffffff",
   47843 => x"ffffff",
   47844 => x"ffffff",
   47845 => x"ffffff",
   47846 => x"ffffff",
   47847 => x"ffffff",
   47848 => x"ffffff",
   47849 => x"ffffff",
   47850 => x"ffffff",
   47851 => x"ffffff",
   47852 => x"ffffff",
   47853 => x"ffffff",
   47854 => x"ffffff",
   47855 => x"ffffff",
   47856 => x"ffffff",
   47857 => x"ffffff",
   47858 => x"ffffff",
   47859 => x"ffffff",
   47860 => x"ffffff",
   47861 => x"ffffff",
   47862 => x"ffffff",
   47863 => x"ffffff",
   47864 => x"ffffff",
   47865 => x"ffffff",
   47866 => x"ffffff",
   47867 => x"ffffff",
   47868 => x"ffffff",
   47869 => x"ffffff",
   47870 => x"ffffff",
   47871 => x"ffffff",
   47872 => x"ffffff",
   47873 => x"ffffff",
   47874 => x"ffffff",
   47875 => x"ffffff",
   47876 => x"ffffff",
   47877 => x"ffffff",
   47878 => x"ffffff",
   47879 => x"ffffff",
   47880 => x"ffffff",
   47881 => x"ffffff",
   47882 => x"ffffff",
   47883 => x"ffffff",
   47884 => x"ffffff",
   47885 => x"ffffff",
   47886 => x"ffffff",
   47887 => x"ffffff",
   47888 => x"ffffff",
   47889 => x"ffffff",
   47890 => x"ffffff",
   47891 => x"ffffff",
   47892 => x"ffffff",
   47893 => x"ffffff",
   47894 => x"ffffff",
   47895 => x"ffffff",
   47896 => x"ffffff",
   47897 => x"ffffff",
   47898 => x"ffffff",
   47899 => x"ffffff",
   47900 => x"ffffff",
   47901 => x"ffffff",
   47902 => x"ffffff",
   47903 => x"ffffff",
   47904 => x"ffffff",
   47905 => x"ffffff",
   47906 => x"ffffff",
   47907 => x"ffffff",
   47908 => x"ffffff",
   47909 => x"fffa95",
   47910 => x"abffff",
   47911 => x"ffffff",
   47912 => x"ffffff",
   47913 => x"ffffff",
   47914 => x"ffffff",
   47915 => x"ffffff",
   47916 => x"ffffff",
   47917 => x"ffffff",
   47918 => x"ffffff",
   47919 => x"ffffff",
   47920 => x"ffffff",
   47921 => x"ffffff",
   47922 => x"ffffff",
   47923 => x"ffffff",
   47924 => x"ffffff",
   47925 => x"ffffff",
   47926 => x"ffffff",
   47927 => x"ffffff",
   47928 => x"ffffff",
   47929 => x"ffffff",
   47930 => x"ffffff",
   47931 => x"ffffff",
   47932 => x"ffffff",
   47933 => x"ffffff",
   47934 => x"ffffff",
   47935 => x"ffffff",
   47936 => x"ffffff",
   47937 => x"ffffff",
   47938 => x"ffffff",
   47939 => x"ffffff",
   47940 => x"ffffff",
   47941 => x"ffffff",
   47942 => x"ffffff",
   47943 => x"ffffff",
   47944 => x"ffffff",
   47945 => x"ffffff",
   47946 => x"ffffff",
   47947 => x"ffffff",
   47948 => x"ffffff",
   47949 => x"ffffff",
   47950 => x"ffffff",
   47951 => x"ffffff",
   47952 => x"ffffff",
   47953 => x"ffffff",
   47954 => x"ffffff",
   47955 => x"ffffff",
   47956 => x"ffffff",
   47957 => x"ffffff",
   47958 => x"ffffff",
   47959 => x"ffffff",
   47960 => x"ffffff",
   47961 => x"ffffff",
   47962 => x"ffffff",
   47963 => x"ffffff",
   47964 => x"ffffff",
   47965 => x"ffffff",
   47966 => x"ffffff",
   47967 => x"ffffff",
   47968 => x"ffffff",
   47969 => x"ffffff",
   47970 => x"ffffff",
   47971 => x"ffffff",
   47972 => x"ffffff",
   47973 => x"ffffff",
   47974 => x"ffffff",
   47975 => x"ffffff",
   47976 => x"ffffff",
   47977 => x"ffffff",
   47978 => x"ffffff",
   47979 => x"ffffff",
   47980 => x"ffffff",
   47981 => x"ffffff",
   47982 => x"ffffff",
   47983 => x"ffffff",
   47984 => x"ffffff",
   47985 => x"ffffff",
   47986 => x"ffffff",
   47987 => x"ffffff",
   47988 => x"ffffff",
   47989 => x"ffffff",
   47990 => x"ffffff",
   47991 => x"ffffff",
   47992 => x"ffffff",
   47993 => x"ffffff",
   47994 => x"ffffff",
   47995 => x"ffffff",
   47996 => x"ffffff",
   47997 => x"ffffff",
   47998 => x"ffffff",
   47999 => x"ffffff",
   48000 => x"ffffff",
   48001 => x"ffffff",
   48002 => x"ffffff",
   48003 => x"ffffff",
   48004 => x"ffffff",
   48005 => x"ffffff",
   48006 => x"ffffff",
   48007 => x"ffffff",
   48008 => x"ffffff",
   48009 => x"ffffff",
   48010 => x"ffffff",
   48011 => x"ffffff",
   48012 => x"ffffff",
   48013 => x"ffffff",
   48014 => x"ffffff",
   48015 => x"ffffff",
   48016 => x"ffffff",
   48017 => x"ffffff",
   48018 => x"ffffff",
   48019 => x"ffffff",
   48020 => x"ffffff",
   48021 => x"ffffff",
   48022 => x"ffffff",
   48023 => x"ffffff",
   48024 => x"ffffff",
   48025 => x"ffffff",
   48026 => x"ffffff",
   48027 => x"ffffff",
   48028 => x"ffffff",
   48029 => x"ffffff",
   48030 => x"ffffff",
   48031 => x"ffffff",
   48032 => x"ffffff",
   48033 => x"ffffff",
   48034 => x"ffffff",
   48035 => x"ffffff",
   48036 => x"ffffff",
   48037 => x"ffffff",
   48038 => x"ffffff",
   48039 => x"ffffff",
   48040 => x"ffffff",
   48041 => x"ffffff",
   48042 => x"ffffff",
   48043 => x"ffffff",
   48044 => x"ffffff",
   48045 => x"ffffff",
   48046 => x"ffffff",
   48047 => x"ffffff",
   48048 => x"ffffff",
   48049 => x"ffffff",
   48050 => x"ffffff",
   48051 => x"ffffff",
   48052 => x"ffffff",
   48053 => x"ffffff",
   48054 => x"ffffff",
   48055 => x"ffffff",
   48056 => x"ffffff",
   48057 => x"ffffff",
   48058 => x"ffffff",
   48059 => x"ffffff",
   48060 => x"ffffff",
   48061 => x"ffffff",
   48062 => x"ffffff",
   48063 => x"ffffff",
   48064 => x"ffffff",
   48065 => x"ffffff",
   48066 => x"ffffff",
   48067 => x"ffffff",
   48068 => x"ffffff",
   48069 => x"fffa95",
   48070 => x"abffff",
   48071 => x"ffffff",
   48072 => x"ffffff",
   48073 => x"ffffff",
   48074 => x"ffffff",
   48075 => x"ffffff",
   48076 => x"ffffff",
   48077 => x"ffffff",
   48078 => x"ffffff",
   48079 => x"ffffff",
   48080 => x"ffffff",
   48081 => x"ffffff",
   48082 => x"ffffff",
   48083 => x"ffffff",
   48084 => x"ffffff",
   48085 => x"ffffff",
   48086 => x"ffffff",
   48087 => x"ffffff",
   48088 => x"ffffff",
   48089 => x"ffffff",
   48090 => x"ffffff",
   48091 => x"ffffff",
   48092 => x"ffffff",
   48093 => x"ffffff",
   48094 => x"ffffff",
   48095 => x"ffffff",
   48096 => x"ffffff",
   48097 => x"ffffff",
   48098 => x"ffffff",
   48099 => x"ffffff",
   48100 => x"ffffff",
   48101 => x"ffffff",
   48102 => x"ffffff",
   48103 => x"ffffff",
   48104 => x"ffffff",
   48105 => x"ffffff",
   48106 => x"ffffff",
   48107 => x"ffffff",
   48108 => x"ffffff",
   48109 => x"ffffff",
   48110 => x"ffffff",
   48111 => x"ffffff",
   48112 => x"ffffff",
   48113 => x"ffffff",
   48114 => x"ffffff",
   48115 => x"ffffff",
   48116 => x"ffffff",
   48117 => x"ffffff",
   48118 => x"ffffff",
   48119 => x"ffffff",
   48120 => x"ffffff",
   48121 => x"ffffff",
   48122 => x"ffffff",
   48123 => x"ffffff",
   48124 => x"ffffff",
   48125 => x"ffffff",
   48126 => x"ffffff",
   48127 => x"ffffff",
   48128 => x"ffffff",
   48129 => x"ffffff",
   48130 => x"ffffff",
   48131 => x"ffffff",
   48132 => x"ffffff",
   48133 => x"ffffff",
   48134 => x"ffffff",
   48135 => x"ffffff",
   48136 => x"ffffff",
   48137 => x"ffffff",
   48138 => x"ffffff",
   48139 => x"ffffff",
   48140 => x"ffffff",
   48141 => x"ffffff",
   48142 => x"ffffff",
   48143 => x"ffffff",
   48144 => x"ffffff",
   48145 => x"ffffff",
   48146 => x"ffffff",
   48147 => x"ffffff",
   48148 => x"ffffff",
   48149 => x"ffffff",
   48150 => x"ffffff",
   48151 => x"ffffff",
   48152 => x"ffffff",
   48153 => x"ffffff",
   48154 => x"ffffff",
   48155 => x"ffffff",
   48156 => x"ffffff",
   48157 => x"ffffff",
   48158 => x"ffffff",
   48159 => x"ffffff",
   48160 => x"ffffff",
   48161 => x"ffffff",
   48162 => x"ffffff",
   48163 => x"ffffff",
   48164 => x"ffffff",
   48165 => x"ffffff",
   48166 => x"ffffff",
   48167 => x"ffffff",
   48168 => x"ffffff",
   48169 => x"ffffff",
   48170 => x"ffffff",
   48171 => x"ffffff",
   48172 => x"ffffff",
   48173 => x"ffffff",
   48174 => x"ffffff",
   48175 => x"ffffff",
   48176 => x"ffffff",
   48177 => x"ffffff",
   48178 => x"ffffff",
   48179 => x"ffffff",
   48180 => x"ffffff",
   48181 => x"ffffff",
   48182 => x"ffffff",
   48183 => x"ffffff",
   48184 => x"ffffff",
   48185 => x"ffffff",
   48186 => x"ffffff",
   48187 => x"ffffff",
   48188 => x"ffffff",
   48189 => x"ffffff",
   48190 => x"ffffff",
   48191 => x"ffffff",
   48192 => x"ffffff",
   48193 => x"ffffff",
   48194 => x"ffffff",
   48195 => x"ffffff",
   48196 => x"ffffff",
   48197 => x"ffffff",
   48198 => x"ffffff",
   48199 => x"ffffff",
   48200 => x"ffffff",
   48201 => x"ffffff",
   48202 => x"ffffff",
   48203 => x"ffffff",
   48204 => x"ffffff",
   48205 => x"ffffff",
   48206 => x"ffffff",
   48207 => x"ffffff",
   48208 => x"ffffff",
   48209 => x"ffffff",
   48210 => x"ffffff",
   48211 => x"ffffff",
   48212 => x"ffffff",
   48213 => x"ffffff",
   48214 => x"ffffff",
   48215 => x"ffffff",
   48216 => x"ffffff",
   48217 => x"ffffff",
   48218 => x"ffffff",
   48219 => x"ffffff",
   48220 => x"ffffff",
   48221 => x"ffffff",
   48222 => x"ffffff",
   48223 => x"ffffff",
   48224 => x"ffffff",
   48225 => x"ffffff",
   48226 => x"ffffff",
   48227 => x"ffffff",
   48228 => x"ffffff",
   48229 => x"fffa95",
   48230 => x"abffff",
   48231 => x"ffffff",
   48232 => x"ffffff",
   48233 => x"ffffff",
   48234 => x"ffffff",
   48235 => x"ffffff",
   48236 => x"ffffff",
   48237 => x"ffffff",
   48238 => x"ffffff",
   48239 => x"ffffff",
   48240 => x"ffffff",
   48241 => x"ffffff",
   48242 => x"ffffff",
   48243 => x"ffffff",
   48244 => x"ffffff",
   48245 => x"ffffff",
   48246 => x"ffffff",
   48247 => x"ffffff",
   48248 => x"ffffff",
   48249 => x"ffffff",
   48250 => x"ffffff",
   48251 => x"ffffff",
   48252 => x"ffffff",
   48253 => x"ffffff",
   48254 => x"ffffff",
   48255 => x"ffffff",
   48256 => x"ffffff",
   48257 => x"ffffff",
   48258 => x"ffffff",
   48259 => x"ffffff",
   48260 => x"ffffff",
   48261 => x"ffffff",
   48262 => x"ffffff",
   48263 => x"ffffff",
   48264 => x"ffffff",
   48265 => x"ffffff",
   48266 => x"ffffff",
   48267 => x"ffffff",
   48268 => x"ffffff",
   48269 => x"ffffff",
   48270 => x"ffffff",
   48271 => x"ffffff",
   48272 => x"ffffff",
   48273 => x"ffffff",
   48274 => x"ffffff",
   48275 => x"ffffff",
   48276 => x"ffffff",
   48277 => x"ffffff",
   48278 => x"ffffff",
   48279 => x"ffffff",
   48280 => x"ffffff",
   48281 => x"ffffff",
   48282 => x"ffffff",
   48283 => x"ffffff",
   48284 => x"ffffff",
   48285 => x"ffffff",
   48286 => x"ffffff",
   48287 => x"ffffff",
   48288 => x"ffffff",
   48289 => x"ffffff",
   48290 => x"ffffff",
   48291 => x"ffffff",
   48292 => x"ffffff",
   48293 => x"ffffff",
   48294 => x"ffffff",
   48295 => x"ffffff",
   48296 => x"ffffff",
   48297 => x"ffffff",
   48298 => x"ffffff",
   48299 => x"ffffff",
   48300 => x"ffffff",
   48301 => x"ffffff",
   48302 => x"ffffff",
   48303 => x"ffffff",
   48304 => x"ffffff",
   48305 => x"ffffff",
   48306 => x"ffffff",
   48307 => x"ffffff",
   48308 => x"ffffff",
   48309 => x"ffffff",
   48310 => x"ffffff",
   48311 => x"ffffff",
   48312 => x"ffffff",
   48313 => x"ffffff",
   48314 => x"ffffff",
   48315 => x"ffffff",
   48316 => x"ffffff",
   48317 => x"ffffff",
   48318 => x"ffffff",
   48319 => x"ffffff",
   48320 => x"ffffff",
   48321 => x"ffffff",
   48322 => x"ffffff",
   48323 => x"ffffff",
   48324 => x"ffffff",
   48325 => x"ffffff",
   48326 => x"ffffff",
   48327 => x"ffffff",
   48328 => x"ffffff",
   48329 => x"ffffff",
   48330 => x"ffffff",
   48331 => x"ffffff",
   48332 => x"ffffff",
   48333 => x"ffffff",
   48334 => x"ffffff",
   48335 => x"ffffff",
   48336 => x"ffffff",
   48337 => x"ffffff",
   48338 => x"ffffff",
   48339 => x"ffffff",
   48340 => x"ffffff",
   48341 => x"ffffff",
   48342 => x"ffffff",
   48343 => x"ffffff",
   48344 => x"ffffff",
   48345 => x"ffffff",
   48346 => x"ffffff",
   48347 => x"ffffff",
   48348 => x"ffffff",
   48349 => x"ffffff",
   48350 => x"ffffff",
   48351 => x"ffffff",
   48352 => x"ffffff",
   48353 => x"ffffff",
   48354 => x"ffffff",
   48355 => x"ffffff",
   48356 => x"ffffff",
   48357 => x"ffffff",
   48358 => x"ffffff",
   48359 => x"ffffff",
   48360 => x"ffffff",
   48361 => x"ffffff",
   48362 => x"ffffff",
   48363 => x"ffffff",
   48364 => x"ffffff",
   48365 => x"ffffff",
   48366 => x"ffffff",
   48367 => x"ffffff",
   48368 => x"ffffff",
   48369 => x"ffffff",
   48370 => x"ffffff",
   48371 => x"ffffff",
   48372 => x"ffffff",
   48373 => x"ffffff",
   48374 => x"ffffff",
   48375 => x"ffffff",
   48376 => x"ffffff",
   48377 => x"ffffff",
   48378 => x"ffffff",
   48379 => x"ffffff",
   48380 => x"ffffff",
   48381 => x"ffffff",
   48382 => x"ffffff",
   48383 => x"ffffff",
   48384 => x"ffffff",
   48385 => x"ffffff",
   48386 => x"ffffff",
   48387 => x"ffffff",
   48388 => x"ffffff",
   48389 => x"fffa95",
   48390 => x"abffff",
   48391 => x"ffffff",
   48392 => x"ffffff",
   48393 => x"ffffff",
   48394 => x"ffffff",
   48395 => x"ffffff",
   48396 => x"ffffff",
   48397 => x"ffffff",
   48398 => x"ffffff",
   48399 => x"ffffff",
   48400 => x"ffffff",
   48401 => x"ffffff",
   48402 => x"ffffff",
   48403 => x"ffffff",
   48404 => x"ffffff",
   48405 => x"ffffff",
   48406 => x"ffffff",
   48407 => x"ffffff",
   48408 => x"ffffff",
   48409 => x"ffffff",
   48410 => x"ffffff",
   48411 => x"ffffff",
   48412 => x"ffffff",
   48413 => x"ffffff",
   48414 => x"ffffff",
   48415 => x"ffffff",
   48416 => x"ffffff",
   48417 => x"ffffff",
   48418 => x"ffffff",
   48419 => x"ffffff",
   48420 => x"ffffff",
   48421 => x"ffffff",
   48422 => x"ffffff",
   48423 => x"ffffff",
   48424 => x"ffffff",
   48425 => x"ffffff",
   48426 => x"ffffff",
   48427 => x"ffffff",
   48428 => x"ffffff",
   48429 => x"ffffff",
   48430 => x"ffffff",
   48431 => x"ffffff",
   48432 => x"ffffff",
   48433 => x"ffffff",
   48434 => x"ffffff",
   48435 => x"ffffff",
   48436 => x"ffffff",
   48437 => x"ffffff",
   48438 => x"ffffff",
   48439 => x"ffffff",
   48440 => x"ffffff",
   48441 => x"ffffff",
   48442 => x"ffffff",
   48443 => x"ffffff",
   48444 => x"ffffff",
   48445 => x"ffffff",
   48446 => x"ffffff",
   48447 => x"ffffff",
   48448 => x"ffffff",
   48449 => x"ffffff",
   48450 => x"ffffff",
   48451 => x"ffffff",
   48452 => x"ffffff",
   48453 => x"ffffff",
   48454 => x"ffffff",
   48455 => x"ffffff",
   48456 => x"ffffff",
   48457 => x"ffffff",
   48458 => x"ffffff",
   48459 => x"ffffff",
   48460 => x"ffffff",
   48461 => x"ffffff",
   48462 => x"ffffff",
   48463 => x"ffffff",
   48464 => x"ffffff",
   48465 => x"ffffff",
   48466 => x"ffffff",
   48467 => x"ffffff",
   48468 => x"ffffff",
   48469 => x"ffffff",
   48470 => x"ffffff",
   48471 => x"ffffff",
   48472 => x"ffffff",
   48473 => x"ffffff",
   48474 => x"ffffff",
   48475 => x"ffffff",
   48476 => x"ffffff",
   48477 => x"ffffff",
   48478 => x"ffffff",
   48479 => x"ffffff",
   48480 => x"ffffff",
   48481 => x"ffffff",
   48482 => x"ffffff",
   48483 => x"ffffff",
   48484 => x"ffffff",
   48485 => x"ffffff",
   48486 => x"ffffff",
   48487 => x"ffffff",
   48488 => x"ffffff",
   48489 => x"ffffff",
   48490 => x"ffffff",
   48491 => x"ffffff",
   48492 => x"ffffff",
   48493 => x"ffffff",
   48494 => x"ffffff",
   48495 => x"ffffff",
   48496 => x"ffffff",
   48497 => x"ffffff",
   48498 => x"ffffff",
   48499 => x"ffffff",
   48500 => x"ffffff",
   48501 => x"ffffff",
   48502 => x"ffffff",
   48503 => x"ffffff",
   48504 => x"ffffff",
   48505 => x"ffffff",
   48506 => x"ffffff",
   48507 => x"ffffff",
   48508 => x"ffffff",
   48509 => x"ffffff",
   48510 => x"ffffff",
   48511 => x"ffffff",
   48512 => x"ffffff",
   48513 => x"ffffff",
   48514 => x"ffffff",
   48515 => x"ffffff",
   48516 => x"ffffff",
   48517 => x"ffffff",
   48518 => x"ffffff",
   48519 => x"ffffff",
   48520 => x"ffffff",
   48521 => x"ffffff",
   48522 => x"ffffff",
   48523 => x"ffffff",
   48524 => x"ffffff",
   48525 => x"ffffff",
   48526 => x"ffffff",
   48527 => x"ffffff",
   48528 => x"ffffff",
   48529 => x"ffffff",
   48530 => x"ffffff",
   48531 => x"ffffff",
   48532 => x"ffffff",
   48533 => x"ffffff",
   48534 => x"ffffff",
   48535 => x"ffffff",
   48536 => x"ffffff",
   48537 => x"ffffff",
   48538 => x"ffffff",
   48539 => x"ffffff",
   48540 => x"ffffff",
   48541 => x"ffffff",
   48542 => x"ffffff",
   48543 => x"ffffff",
   48544 => x"ffffff",
   48545 => x"ffffff",
   48546 => x"ffffff",
   48547 => x"ffffff",
   48548 => x"ffffff",
   48549 => x"fffa95",
   48550 => x"abffff",
   48551 => x"ffffff",
   48552 => x"ffffff",
   48553 => x"ffffff",
   48554 => x"ffffff",
   48555 => x"ffffff",
   48556 => x"ffffff",
   48557 => x"ffffff",
   48558 => x"ffffff",
   48559 => x"ffffff",
   48560 => x"ffffff",
   48561 => x"ffffff",
   48562 => x"ffffff",
   48563 => x"ffffff",
   48564 => x"ffffff",
   48565 => x"ffffff",
   48566 => x"ffffff",
   48567 => x"ffffff",
   48568 => x"ffffff",
   48569 => x"ffffff",
   48570 => x"ffffff",
   48571 => x"ffffff",
   48572 => x"ffffff",
   48573 => x"ffffff",
   48574 => x"ffffff",
   48575 => x"ffffff",
   48576 => x"ffffff",
   48577 => x"ffffff",
   48578 => x"ffffff",
   48579 => x"ffffff",
   48580 => x"ffffff",
   48581 => x"ffffff",
   48582 => x"ffffff",
   48583 => x"ffffff",
   48584 => x"ffffff",
   48585 => x"ffffff",
   48586 => x"ffffff",
   48587 => x"ffffff",
   48588 => x"ffffff",
   48589 => x"ffffff",
   48590 => x"ffffff",
   48591 => x"ffffff",
   48592 => x"ffffff",
   48593 => x"ffffff",
   48594 => x"ffffff",
   48595 => x"ffffff",
   48596 => x"ffffff",
   48597 => x"ffffff",
   48598 => x"ffffff",
   48599 => x"ffffff",
   48600 => x"ffffff",
   48601 => x"ffffff",
   48602 => x"ffffff",
   48603 => x"ffffff",
   48604 => x"ffffff",
   48605 => x"ffffff",
   48606 => x"ffffff",
   48607 => x"ffffff",
   48608 => x"ffffff",
   48609 => x"ffffff",
   48610 => x"ffffff",
   48611 => x"ffffff",
   48612 => x"ffffff",
   48613 => x"ffffff",
   48614 => x"ffffff",
   48615 => x"ffffff",
   48616 => x"ffffff",
   48617 => x"ffffff",
   48618 => x"ffffff",
   48619 => x"ffffff",
   48620 => x"ffffff",
   48621 => x"ffffff",
   48622 => x"ffffff",
   48623 => x"ffffff",
   48624 => x"ffffff",
   48625 => x"ffffff",
   48626 => x"ffffff",
   48627 => x"ffffff",
   48628 => x"ffffff",
   48629 => x"ffffff",
   48630 => x"ffffff",
   48631 => x"ffffff",
   48632 => x"ffffff",
   48633 => x"ffffff",
   48634 => x"ffffff",
   48635 => x"ffffff",
   48636 => x"ffffff",
   48637 => x"ffffff",
   48638 => x"ffffff",
   48639 => x"ffffff",
   48640 => x"ffffff",
   48641 => x"ffffff",
   48642 => x"ffffff",
   48643 => x"ffffff",
   48644 => x"ffffff",
   48645 => x"ffffff",
   48646 => x"ffffff",
   48647 => x"ffffff",
   48648 => x"ffffff",
   48649 => x"ffffff",
   48650 => x"ffffff",
   48651 => x"ffffff",
   48652 => x"ffffff",
   48653 => x"ffffff",
   48654 => x"ffffff",
   48655 => x"ffffff",
   48656 => x"ffffff",
   48657 => x"ffffff",
   48658 => x"ffffff",
   48659 => x"ffffff",
   48660 => x"ffffff",
   48661 => x"ffffff",
   48662 => x"ffffff",
   48663 => x"ffffff",
   48664 => x"ffffff",
   48665 => x"ffffff",
   48666 => x"ffffff",
   48667 => x"ffffff",
   48668 => x"ffffff",
   48669 => x"ffffff",
   48670 => x"ffffff",
   48671 => x"ffffff",
   48672 => x"ffffff",
   48673 => x"ffffff",
   48674 => x"ffffff",
   48675 => x"ffffff",
   48676 => x"ffffff",
   48677 => x"ffffff",
   48678 => x"ffffff",
   48679 => x"ffffff",
   48680 => x"ffffff",
   48681 => x"ffffff",
   48682 => x"ffffff",
   48683 => x"ffffff",
   48684 => x"ffffff",
   48685 => x"ffffff",
   48686 => x"ffffff",
   48687 => x"ffffff",
   48688 => x"ffffff",
   48689 => x"ffffff",
   48690 => x"ffffff",
   48691 => x"ffffff",
   48692 => x"ffffff",
   48693 => x"ffffff",
   48694 => x"ffffff",
   48695 => x"ffffff",
   48696 => x"ffffff",
   48697 => x"ffffff",
   48698 => x"ffffff",
   48699 => x"ffffff",
   48700 => x"ffffff",
   48701 => x"ffffff",
   48702 => x"ffffff",
   48703 => x"ffffff",
   48704 => x"ffffff",
   48705 => x"ffffff",
   48706 => x"ffffff",
   48707 => x"ffffff",
   48708 => x"ffffff",
   48709 => x"fffa95",
   48710 => x"abffff",
   48711 => x"ffffff",
   48712 => x"ffffff",
   48713 => x"ffffff",
   48714 => x"ffffff",
   48715 => x"ffffff",
   48716 => x"ffffff",
   48717 => x"ffffff",
   48718 => x"ffffff",
   48719 => x"ffffff",
   48720 => x"ffffff",
   48721 => x"ffffff",
   48722 => x"ffffff",
   48723 => x"ffffff",
   48724 => x"ffffff",
   48725 => x"ffffff",
   48726 => x"ffffff",
   48727 => x"ffffff",
   48728 => x"ffffff",
   48729 => x"ffffff",
   48730 => x"ffffff",
   48731 => x"ffffff",
   48732 => x"ffffff",
   48733 => x"ffffff",
   48734 => x"ffffff",
   48735 => x"ffffff",
   48736 => x"ffffff",
   48737 => x"ffffff",
   48738 => x"ffffff",
   48739 => x"ffffff",
   48740 => x"ffffff",
   48741 => x"ffffff",
   48742 => x"ffffff",
   48743 => x"ffffff",
   48744 => x"ffffff",
   48745 => x"ffffff",
   48746 => x"ffffff",
   48747 => x"ffffff",
   48748 => x"ffffff",
   48749 => x"ffffff",
   48750 => x"ffffff",
   48751 => x"ffffff",
   48752 => x"ffffff",
   48753 => x"ffffff",
   48754 => x"ffffff",
   48755 => x"ffffff",
   48756 => x"ffffff",
   48757 => x"ffffff",
   48758 => x"ffffff",
   48759 => x"ffffff",
   48760 => x"ffffff",
   48761 => x"ffffff",
   48762 => x"ffffff",
   48763 => x"ffffff",
   48764 => x"ffffff",
   48765 => x"ffffff",
   48766 => x"ffffff",
   48767 => x"ffffff",
   48768 => x"ffffff",
   48769 => x"ffffff",
   48770 => x"ffffff",
   48771 => x"ffffff",
   48772 => x"ffffff",
   48773 => x"ffffff",
   48774 => x"ffffff",
   48775 => x"ffffff",
   48776 => x"ffffff",
   48777 => x"ffffff",
   48778 => x"ffffff",
   48779 => x"ffffff",
   48780 => x"ffffff",
   48781 => x"ffffff",
   48782 => x"ffffff",
   48783 => x"ffffff",
   48784 => x"ffffff",
   48785 => x"ffffff",
   48786 => x"ffffff",
   48787 => x"ffffff",
   48788 => x"ffffff",
   48789 => x"ffffff",
   48790 => x"ffffff",
   48791 => x"ffffff",
   48792 => x"ffffff",
   48793 => x"ffffff",
   48794 => x"ffffff",
   48795 => x"ffffff",
   48796 => x"ffffff",
   48797 => x"ffffff",
   48798 => x"ffffff",
   48799 => x"ffffff",
   48800 => x"ffffff",
   48801 => x"ffffff",
   48802 => x"ffffff",
   48803 => x"ffffff",
   48804 => x"ffffff",
   48805 => x"ffffff",
   48806 => x"ffffff",
   48807 => x"ffffff",
   48808 => x"ffffff",
   48809 => x"ffffff",
   48810 => x"ffffff",
   48811 => x"ffffff",
   48812 => x"ffffff",
   48813 => x"ffffff",
   48814 => x"ffffff",
   48815 => x"ffffff",
   48816 => x"ffffff",
   48817 => x"ffffff",
   48818 => x"ffffff",
   48819 => x"ffffff",
   48820 => x"ffffff",
   48821 => x"ffffff",
   48822 => x"ffffff",
   48823 => x"ffffff",
   48824 => x"ffffff",
   48825 => x"ffffff",
   48826 => x"ffffff",
   48827 => x"ffffff",
   48828 => x"ffffff",
   48829 => x"ffffff",
   48830 => x"ffffff",
   48831 => x"ffffff",
   48832 => x"ffffff",
   48833 => x"ffffff",
   48834 => x"ffffff",
   48835 => x"ffffff",
   48836 => x"ffffff",
   48837 => x"ffffff",
   48838 => x"ffffff",
   48839 => x"ffffff",
   48840 => x"ffffff",
   48841 => x"ffffff",
   48842 => x"ffffff",
   48843 => x"ffffff",
   48844 => x"ffffff",
   48845 => x"ffffff",
   48846 => x"ffffff",
   48847 => x"ffffff",
   48848 => x"ffffff",
   48849 => x"ffffff",
   48850 => x"ffffff",
   48851 => x"ffffff",
   48852 => x"ffffff",
   48853 => x"ffffff",
   48854 => x"ffffff",
   48855 => x"ffffff",
   48856 => x"ffffff",
   48857 => x"ffffff",
   48858 => x"ffffff",
   48859 => x"ffffff",
   48860 => x"ffffff",
   48861 => x"ffffff",
   48862 => x"ffffff",
   48863 => x"ffffff",
   48864 => x"ffffff",
   48865 => x"ffffff",
   48866 => x"ffffff",
   48867 => x"ffffff",
   48868 => x"ffffff",
   48869 => x"fffa95",
   48870 => x"abffff",
   48871 => x"ffffff",
   48872 => x"ffffff",
   48873 => x"ffffff",
   48874 => x"ffffff",
   48875 => x"ffffff",
   48876 => x"ffffff",
   48877 => x"ffffff",
   48878 => x"ffffff",
   48879 => x"ffffff",
   48880 => x"ffffff",
   48881 => x"ffffff",
   48882 => x"ffffff",
   48883 => x"ffffff",
   48884 => x"ffffff",
   48885 => x"ffffff",
   48886 => x"ffffff",
   48887 => x"ffffff",
   48888 => x"ffffff",
   48889 => x"ffffff",
   48890 => x"ffffff",
   48891 => x"ffffff",
   48892 => x"ffffff",
   48893 => x"ffffff",
   48894 => x"ffffff",
   48895 => x"ffffff",
   48896 => x"ffffff",
   48897 => x"ffffff",
   48898 => x"ffffff",
   48899 => x"ffffff",
   48900 => x"ffffff",
   48901 => x"ffffff",
   48902 => x"ffffff",
   48903 => x"ffffff",
   48904 => x"ffffff",
   48905 => x"ffffff",
   48906 => x"ffffff",
   48907 => x"ffffff",
   48908 => x"ffffff",
   48909 => x"ffffff",
   48910 => x"ffffff",
   48911 => x"ffffff",
   48912 => x"ffffff",
   48913 => x"ffffff",
   48914 => x"ffffff",
   48915 => x"ffffff",
   48916 => x"ffffff",
   48917 => x"ffffff",
   48918 => x"ffffff",
   48919 => x"ffffff",
   48920 => x"ffffff",
   48921 => x"ffffff",
   48922 => x"ffffff",
   48923 => x"ffffff",
   48924 => x"ffffff",
   48925 => x"ffffff",
   48926 => x"ffffff",
   48927 => x"ffffff",
   48928 => x"ffffff",
   48929 => x"ffffff",
   48930 => x"ffffff",
   48931 => x"ffffff",
   48932 => x"ffffff",
   48933 => x"ffffff",
   48934 => x"ffffff",
   48935 => x"ffffff",
   48936 => x"ffffff",
   48937 => x"ffffff",
   48938 => x"ffffff",
   48939 => x"ffffff",
   48940 => x"ffffff",
   48941 => x"ffffff",
   48942 => x"ffffff",
   48943 => x"ffffff",
   48944 => x"ffffff",
   48945 => x"ffffff",
   48946 => x"ffffff",
   48947 => x"ffffff",
   48948 => x"ffffff",
   48949 => x"ffffff",
   48950 => x"ffffff",
   48951 => x"ffffff",
   48952 => x"ffffff",
   48953 => x"ffffff",
   48954 => x"ffffff",
   48955 => x"ffffff",
   48956 => x"ffffff",
   48957 => x"ffffff",
   48958 => x"ffffff",
   48959 => x"ffffff",
   48960 => x"ffffff",
   48961 => x"ffffff",
   48962 => x"ffffff",
   48963 => x"ffffff",
   48964 => x"ffffff",
   48965 => x"ffffff",
   48966 => x"ffffff",
   48967 => x"ffffff",
   48968 => x"ffffff",
   48969 => x"ffffff",
   48970 => x"ffffff",
   48971 => x"ffffff",
   48972 => x"ffffff",
   48973 => x"ffffff",
   48974 => x"ffffff",
   48975 => x"ffffff",
   48976 => x"ffffff",
   48977 => x"ffffff",
   48978 => x"ffffff",
   48979 => x"ffffff",
   48980 => x"ffffff",
   48981 => x"ffffff",
   48982 => x"ffffff",
   48983 => x"ffffff",
   48984 => x"ffffff",
   48985 => x"ffffff",
   48986 => x"ffffff",
   48987 => x"ffffff",
   48988 => x"ffffff",
   48989 => x"ffffff",
   48990 => x"ffffff",
   48991 => x"ffffff",
   48992 => x"ffffff",
   48993 => x"ffffff",
   48994 => x"ffffff",
   48995 => x"ffffff",
   48996 => x"ffffff",
   48997 => x"ffffff",
   48998 => x"ffffff",
   48999 => x"ffffff",
   49000 => x"ffffff",
   49001 => x"ffffff",
   49002 => x"ffffff",
   49003 => x"ffffff",
   49004 => x"ffffff",
   49005 => x"ffffff",
   49006 => x"ffffff",
   49007 => x"ffffff",
   49008 => x"ffffff",
   49009 => x"ffffff",
   49010 => x"ffffff",
   49011 => x"ffffff",
   49012 => x"ffffff",
   49013 => x"ffffff",
   49014 => x"ffffff",
   49015 => x"ffffff",
   49016 => x"ffffff",
   49017 => x"ffffff",
   49018 => x"ffffff",
   49019 => x"ffffff",
   49020 => x"ffffff",
   49021 => x"ffffff",
   49022 => x"ffffff",
   49023 => x"ffffff",
   49024 => x"ffffff",
   49025 => x"ffffff",
   49026 => x"ffffff",
   49027 => x"ffffff",
   49028 => x"ffffff",
   49029 => x"fffa95",
   49030 => x"abffff",
   49031 => x"ffffff",
   49032 => x"ffffff",
   49033 => x"ffffff",
   49034 => x"ffffff",
   49035 => x"ffffff",
   49036 => x"ffffff",
   49037 => x"ffffff",
   49038 => x"ffffff",
   49039 => x"ffffff",
   49040 => x"ffffff",
   49041 => x"ffffff",
   49042 => x"ffffff",
   49043 => x"ffffff",
   49044 => x"ffffff",
   49045 => x"ffffff",
   49046 => x"ffffff",
   49047 => x"ffffff",
   49048 => x"ffffff",
   49049 => x"ffffff",
   49050 => x"ffffff",
   49051 => x"ffffff",
   49052 => x"ffffff",
   49053 => x"ffffff",
   49054 => x"ffffff",
   49055 => x"ffffff",
   49056 => x"ffffff",
   49057 => x"ffffff",
   49058 => x"ffffff",
   49059 => x"ffffff",
   49060 => x"ffffff",
   49061 => x"ffffff",
   49062 => x"ffffff",
   49063 => x"ffffff",
   49064 => x"ffffff",
   49065 => x"ffffff",
   49066 => x"ffffff",
   49067 => x"ffffff",
   49068 => x"ffffff",
   49069 => x"ffffff",
   49070 => x"ffffff",
   49071 => x"ffffff",
   49072 => x"ffffff",
   49073 => x"ffffff",
   49074 => x"ffffff",
   49075 => x"ffffff",
   49076 => x"ffffff",
   49077 => x"ffffff",
   49078 => x"ffffff",
   49079 => x"ffffff",
   49080 => x"ffffff",
   49081 => x"ffffff",
   49082 => x"ffffff",
   49083 => x"ffffff",
   49084 => x"ffffff",
   49085 => x"ffffff",
   49086 => x"ffffff",
   49087 => x"ffffff",
   49088 => x"ffffff",
   49089 => x"ffffff",
   49090 => x"ffffff",
   49091 => x"ffffff",
   49092 => x"ffffff",
   49093 => x"ffffff",
   49094 => x"ffffff",
   49095 => x"ffffff",
   49096 => x"ffffff",
   49097 => x"ffffff",
   49098 => x"ffffff",
   49099 => x"ffffff",
   49100 => x"ffffff",
   49101 => x"ffffff",
   49102 => x"ffffff",
   49103 => x"ffffff",
   49104 => x"ffffff",
   49105 => x"ffffff",
   49106 => x"ffffff",
   49107 => x"ffffff",
   49108 => x"ffffff",
   49109 => x"ffffff",
   49110 => x"ffffff",
   49111 => x"ffffff",
   49112 => x"ffffff",
   49113 => x"ffffff",
   49114 => x"ffffff",
   49115 => x"ffffff",
   49116 => x"ffffff",
   49117 => x"ffffff",
   49118 => x"ffffff",
   49119 => x"ffffff",
   49120 => x"ffffff",
   49121 => x"ffffff",
   49122 => x"ffffff",
   49123 => x"ffffff",
   49124 => x"ffffff",
   49125 => x"ffffff",
   49126 => x"ffffff",
   49127 => x"ffffff",
   49128 => x"ffffff",
   49129 => x"ffffff",
   49130 => x"ffffff",
   49131 => x"ffffff",
   49132 => x"ffffff",
   49133 => x"ffffff",
   49134 => x"ffffff",
   49135 => x"ffffff",
   49136 => x"ffffff",
   49137 => x"ffffff",
   49138 => x"ffffff",
   49139 => x"ffffff",
   49140 => x"ffffff",
   49141 => x"ffffff",
   49142 => x"ffffff",
   49143 => x"ffffff",
   49144 => x"ffffff",
   49145 => x"ffffff",
   49146 => x"ffffff",
   49147 => x"ffffff",
   49148 => x"ffffff",
   49149 => x"ffffff",
   49150 => x"ffffff",
   49151 => x"ffffff",
   49152 => x"ffffff",
   49153 => x"ffffff",
   49154 => x"ffffff",
   49155 => x"ffffff",
   49156 => x"ffffff",
   49157 => x"ffffff",
   49158 => x"ffffff",
   49159 => x"ffffff",
   49160 => x"ffffff",
   49161 => x"ffffff",
   49162 => x"ffffff",
   49163 => x"ffffff",
   49164 => x"ffffff",
   49165 => x"ffffff",
   49166 => x"ffffff",
   49167 => x"ffffff",
   49168 => x"ffffff",
   49169 => x"ffffff",
   49170 => x"ffffff",
   49171 => x"ffffff",
   49172 => x"ffffff",
   49173 => x"ffffff",
   49174 => x"ffffff",
   49175 => x"ffffff",
   49176 => x"ffffff",
   49177 => x"ffffff",
   49178 => x"ffffff",
   49179 => x"ffffff",
   49180 => x"ffffff",
   49181 => x"ffffff",
   49182 => x"ffffff",
   49183 => x"ffffff",
   49184 => x"ffffff",
   49185 => x"ffffff",
   49186 => x"ffffff",
   49187 => x"ffffff",
   49188 => x"ffffff",
   49189 => x"fffa95",
   49190 => x"abffff",
   49191 => x"ffffff",
   49192 => x"ffffff",
   49193 => x"ffffff",
   49194 => x"ffffff",
   49195 => x"ffffff",
   49196 => x"ffffff",
   49197 => x"ffffff",
   49198 => x"ffffff",
   49199 => x"ffffff",
   49200 => x"ffffff",
   49201 => x"ffffff",
   49202 => x"ffffff",
   49203 => x"ffffff",
   49204 => x"ffffff",
   49205 => x"ffffff",
   49206 => x"ffffff",
   49207 => x"ffffff",
   49208 => x"ffffff",
   49209 => x"ffffff",
   49210 => x"ffffff",
   49211 => x"ffffff",
   49212 => x"ffffff",
   49213 => x"ffffff",
   49214 => x"ffffff",
   49215 => x"ffffff",
   49216 => x"ffffff",
   49217 => x"ffffff",
   49218 => x"ffffff",
   49219 => x"ffffff",
   49220 => x"ffffff",
   49221 => x"ffffff",
   49222 => x"ffffff",
   49223 => x"ffffff",
   49224 => x"ffffff",
   49225 => x"ffffff",
   49226 => x"ffffff",
   49227 => x"ffffff",
   49228 => x"ffffff",
   49229 => x"ffffff",
   49230 => x"ffffff",
   49231 => x"ffffff",
   49232 => x"ffffff",
   49233 => x"ffffff",
   49234 => x"ffffff",
   49235 => x"ffffff",
   49236 => x"ffffff",
   49237 => x"ffffff",
   49238 => x"ffffff",
   49239 => x"ffffff",
   49240 => x"ffffff",
   49241 => x"ffffff",
   49242 => x"ffffff",
   49243 => x"ffffff",
   49244 => x"ffffff",
   49245 => x"ffffff",
   49246 => x"ffffff",
   49247 => x"ffffff",
   49248 => x"ffffff",
   49249 => x"ffffff",
   49250 => x"ffffff",
   49251 => x"ffffff",
   49252 => x"ffffff",
   49253 => x"ffffff",
   49254 => x"ffffff",
   49255 => x"ffffff",
   49256 => x"ffffff",
   49257 => x"ffffff",
   49258 => x"ffffff",
   49259 => x"ffffff",
   49260 => x"ffffff",
   49261 => x"ffffff",
   49262 => x"ffffff",
   49263 => x"ffffff",
   49264 => x"ffffff",
   49265 => x"ffffff",
   49266 => x"ffffff",
   49267 => x"ffffff",
   49268 => x"ffffff",
   49269 => x"ffffff",
   49270 => x"ffffff",
   49271 => x"ffffff",
   49272 => x"ffffff",
   49273 => x"ffffff",
   49274 => x"ffffff",
   49275 => x"ffffff",
   49276 => x"ffffff",
   49277 => x"ffffff",
   49278 => x"ffffff",
   49279 => x"ffffff",
   49280 => x"ffffff",
   49281 => x"ffffff",
   49282 => x"ffffff",
   49283 => x"ffffff",
   49284 => x"ffffff",
   49285 => x"ffffff",
   49286 => x"ffffff",
   49287 => x"ffffff",
   49288 => x"ffffff",
   49289 => x"ffffff",
   49290 => x"ffffff",
   49291 => x"ffffff",
   49292 => x"ffffff",
   49293 => x"ffffff",
   49294 => x"ffffff",
   49295 => x"ffffff",
   49296 => x"ffffff",
   49297 => x"ffffff",
   49298 => x"ffffff",
   49299 => x"ffffff",
   49300 => x"ffffff",
   49301 => x"ffffff",
   49302 => x"ffffff",
   49303 => x"ffffff",
   49304 => x"ffffff",
   49305 => x"ffffff",
   49306 => x"ffffff",
   49307 => x"ffffff",
   49308 => x"ffffff",
   49309 => x"ffffff",
   49310 => x"ffffff",
   49311 => x"ffffff",
   49312 => x"ffffff",
   49313 => x"ffffff",
   49314 => x"ffffff",
   49315 => x"ffffff",
   49316 => x"ffffff",
   49317 => x"ffffff",
   49318 => x"ffffff",
   49319 => x"ffffff",
   49320 => x"ffffff",
   49321 => x"ffffff",
   49322 => x"ffffff",
   49323 => x"ffffff",
   49324 => x"ffffff",
   49325 => x"ffffff",
   49326 => x"ffffff",
   49327 => x"ffffff",
   49328 => x"ffffff",
   49329 => x"ffffff",
   49330 => x"ffffff",
   49331 => x"ffffff",
   49332 => x"ffffff",
   49333 => x"ffffff",
   49334 => x"ffffff",
   49335 => x"ffffff",
   49336 => x"ffffff",
   49337 => x"ffffff",
   49338 => x"ffffff",
   49339 => x"ffffff",
   49340 => x"ffffff",
   49341 => x"ffffff",
   49342 => x"ffffff",
   49343 => x"ffffff",
   49344 => x"ffffff",
   49345 => x"ffffff",
   49346 => x"ffffff",
   49347 => x"ffffff",
   49348 => x"ffffff",
   49349 => x"fffa95",
   49350 => x"abffff",
   49351 => x"ffffff",
   49352 => x"ffffff",
   49353 => x"ffffff",
   49354 => x"ffffff",
   49355 => x"ffffff",
   49356 => x"ffffff",
   49357 => x"ffffff",
   49358 => x"ffffff",
   49359 => x"ffffff",
   49360 => x"ffffff",
   49361 => x"ffffff",
   49362 => x"ffffff",
   49363 => x"ffffff",
   49364 => x"ffffff",
   49365 => x"ffffff",
   49366 => x"ffffff",
   49367 => x"ffffff",
   49368 => x"ffffff",
   49369 => x"ffffff",
   49370 => x"ffffff",
   49371 => x"ffffff",
   49372 => x"ffffff",
   49373 => x"ffffff",
   49374 => x"ffffff",
   49375 => x"ffffff",
   49376 => x"ffffff",
   49377 => x"ffffff",
   49378 => x"ffffff",
   49379 => x"ffffff",
   49380 => x"ffffff",
   49381 => x"ffffff",
   49382 => x"ffffff",
   49383 => x"ffffff",
   49384 => x"ffffff",
   49385 => x"ffffff",
   49386 => x"ffffff",
   49387 => x"ffffff",
   49388 => x"ffffff",
   49389 => x"ffffff",
   49390 => x"ffffff",
   49391 => x"ffffff",
   49392 => x"ffffff",
   49393 => x"ffffff",
   49394 => x"ffffff",
   49395 => x"ffffff",
   49396 => x"ffffff",
   49397 => x"ffffff",
   49398 => x"ffffff",
   49399 => x"ffffff",
   49400 => x"ffffff",
   49401 => x"ffffff",
   49402 => x"ffffff",
   49403 => x"ffffff",
   49404 => x"ffffff",
   49405 => x"ffffff",
   49406 => x"ffffff",
   49407 => x"ffffff",
   49408 => x"ffffff",
   49409 => x"ffffff",
   49410 => x"ffffff",
   49411 => x"ffffff",
   49412 => x"ffffff",
   49413 => x"ffffff",
   49414 => x"ffffff",
   49415 => x"ffffff",
   49416 => x"ffffff",
   49417 => x"ffffff",
   49418 => x"ffffff",
   49419 => x"ffffff",
   49420 => x"ffffff",
   49421 => x"ffffff",
   49422 => x"ffffff",
   49423 => x"ffffff",
   49424 => x"ffffff",
   49425 => x"ffffff",
   49426 => x"ffffff",
   49427 => x"ffffff",
   49428 => x"ffffff",
   49429 => x"feafff",
   49430 => x"ffffff",
   49431 => x"ffffff",
   49432 => x"ffffff",
   49433 => x"ffffff",
   49434 => x"ffffff",
   49435 => x"ffffff",
   49436 => x"ffffff",
   49437 => x"ffffff",
   49438 => x"ffffff",
   49439 => x"ffffff",
   49440 => x"ffffff",
   49441 => x"ffffff",
   49442 => x"ffffff",
   49443 => x"ffffff",
   49444 => x"ffffff",
   49445 => x"ffffff",
   49446 => x"ffffff",
   49447 => x"ffffff",
   49448 => x"ffffff",
   49449 => x"ffffff",
   49450 => x"ffffff",
   49451 => x"ffffff",
   49452 => x"ffffff",
   49453 => x"ffffff",
   49454 => x"ffffff",
   49455 => x"ffffff",
   49456 => x"ffffff",
   49457 => x"ffffff",
   49458 => x"ffffff",
   49459 => x"ffffff",
   49460 => x"ffffff",
   49461 => x"ffffff",
   49462 => x"ffffff",
   49463 => x"ffffff",
   49464 => x"ffffff",
   49465 => x"ffffff",
   49466 => x"ffffff",
   49467 => x"ffffff",
   49468 => x"ffffff",
   49469 => x"ffffff",
   49470 => x"ffffff",
   49471 => x"ffffff",
   49472 => x"ffffff",
   49473 => x"ffffff",
   49474 => x"ffffff",
   49475 => x"ffffff",
   49476 => x"ffffff",
   49477 => x"ffffff",
   49478 => x"ffffff",
   49479 => x"ffffff",
   49480 => x"ffffff",
   49481 => x"ffffff",
   49482 => x"ffffff",
   49483 => x"ffffff",
   49484 => x"ffffff",
   49485 => x"ffffff",
   49486 => x"ffffff",
   49487 => x"ffffff",
   49488 => x"ffffff",
   49489 => x"ffffff",
   49490 => x"ffffff",
   49491 => x"ffffff",
   49492 => x"ffffff",
   49493 => x"ffffff",
   49494 => x"ffffff",
   49495 => x"ffffff",
   49496 => x"ffffff",
   49497 => x"ffffff",
   49498 => x"ffffff",
   49499 => x"ffffff",
   49500 => x"ffffff",
   49501 => x"ffffff",
   49502 => x"ffffff",
   49503 => x"ffffff",
   49504 => x"ffffff",
   49505 => x"ffffff",
   49506 => x"ffffff",
   49507 => x"ffffff",
   49508 => x"ffffff",
   49509 => x"fffa95",
   49510 => x"abffff",
   49511 => x"ffffff",
   49512 => x"ffffff",
   49513 => x"ffffff",
   49514 => x"ffffff",
   49515 => x"ffffff",
   49516 => x"ffffff",
   49517 => x"ffffff",
   49518 => x"ffffff",
   49519 => x"ffffff",
   49520 => x"ffffff",
   49521 => x"fffad7",
   49522 => x"5d75d7",
   49523 => x"5d75d7",
   49524 => x"5d75d7",
   49525 => x"5d75d7",
   49526 => x"5d75d7",
   49527 => x"5d75d7",
   49528 => x"5d75d7",
   49529 => x"5d75d7",
   49530 => x"5d75d7",
   49531 => x"5d75d7",
   49532 => x"5d75d7",
   49533 => x"5d75d7",
   49534 => x"5d75d7",
   49535 => x"5d75d7",
   49536 => x"5d75d6",
   49537 => x"596596",
   49538 => x"596596",
   49539 => x"596596",
   49540 => x"596596",
   49541 => x"596596",
   49542 => x"596596",
   49543 => x"596596",
   49544 => x"596596",
   49545 => x"596596",
   49546 => x"596596",
   49547 => x"596596",
   49548 => x"596596",
   49549 => x"596596",
   49550 => x"596596",
   49551 => x"596596",
   49552 => x"596596",
   49553 => x"596596",
   49554 => x"596596",
   49555 => x"596596",
   49556 => x"596596",
   49557 => x"596596",
   49558 => x"596596",
   49559 => x"596596",
   49560 => x"596596",
   49561 => x"596596",
   49562 => x"596596",
   49563 => x"596596",
   49564 => x"596596",
   49565 => x"596596",
   49566 => x"596596",
   49567 => x"595555",
   49568 => x"555555",
   49569 => x"555555",
   49570 => x"555555",
   49571 => x"555555",
   49572 => x"555555",
   49573 => x"555555",
   49574 => x"555555",
   49575 => x"555555",
   49576 => x"555555",
   49577 => x"555555",
   49578 => x"555555",
   49579 => x"555555",
   49580 => x"555555",
   49581 => x"555555",
   49582 => x"555555",
   49583 => x"555555",
   49584 => x"555555",
   49585 => x"555555",
   49586 => x"555555",
   49587 => x"555555",
   49588 => x"555555",
   49589 => x"555abf",
   49590 => x"ffffff",
   49591 => x"ffffff",
   49592 => x"ffffff",
   49593 => x"ffffff",
   49594 => x"ffffff",
   49595 => x"ffffff",
   49596 => x"ffffff",
   49597 => x"ffffff",
   49598 => x"ffffff",
   49599 => x"ffffff",
   49600 => x"ffffff",
   49601 => x"ffffff",
   49602 => x"ffffff",
   49603 => x"ffffff",
   49604 => x"ffffff",
   49605 => x"ffffff",
   49606 => x"ffffff",
   49607 => x"ffffff",
   49608 => x"ffffff",
   49609 => x"ffffff",
   49610 => x"ffffff",
   49611 => x"ffffff",
   49612 => x"ffffff",
   49613 => x"ffffff",
   49614 => x"ffffff",
   49615 => x"ffffff",
   49616 => x"ffffff",
   49617 => x"ffffff",
   49618 => x"ffffff",
   49619 => x"ffffff",
   49620 => x"ffffff",
   49621 => x"ffffff",
   49622 => x"ffffff",
   49623 => x"ffffff",
   49624 => x"ffffff",
   49625 => x"ffffff",
   49626 => x"ffffff",
   49627 => x"ffffff",
   49628 => x"ffffff",
   49629 => x"ffffff",
   49630 => x"ffffff",
   49631 => x"ffffff",
   49632 => x"ffffff",
   49633 => x"ffffff",
   49634 => x"ffffff",
   49635 => x"ffffff",
   49636 => x"ffffff",
   49637 => x"ffffff",
   49638 => x"ffffff",
   49639 => x"ffffff",
   49640 => x"ffffff",
   49641 => x"ffffff",
   49642 => x"ffffff",
   49643 => x"ffffff",
   49644 => x"ffffff",
   49645 => x"ffffff",
   49646 => x"ffffff",
   49647 => x"ffffff",
   49648 => x"ffffff",
   49649 => x"ffffff",
   49650 => x"ffffff",
   49651 => x"ffffff",
   49652 => x"ffffff",
   49653 => x"ffffff",
   49654 => x"ffffff",
   49655 => x"ffffff",
   49656 => x"ffffff",
   49657 => x"ffffff",
   49658 => x"ffffff",
   49659 => x"ffffff",
   49660 => x"ffffff",
   49661 => x"ffffff",
   49662 => x"ffffff",
   49663 => x"ffffff",
   49664 => x"ffffff",
   49665 => x"ffffff",
   49666 => x"ffffff",
   49667 => x"ffffff",
   49668 => x"ffffff",
   49669 => x"fffa95",
   49670 => x"abffff",
   49671 => x"ffffff",
   49672 => x"ffffff",
   49673 => x"ffffff",
   49674 => x"ffffff",
   49675 => x"ffffff",
   49676 => x"ffffff",
   49677 => x"ffffff",
   49678 => x"ffffff",
   49679 => x"ffffff",
   49680 => x"ffffff",
   49681 => x"fffac3",
   49682 => x"0c30c3",
   49683 => x"0c30c3",
   49684 => x"0c30c3",
   49685 => x"0c30c3",
   49686 => x"0c30c3",
   49687 => x"0c30c3",
   49688 => x"0c30c3",
   49689 => x"0c30c3",
   49690 => x"0c30c3",
   49691 => x"0c30c3",
   49692 => x"0c30c3",
   49693 => x"082082",
   49694 => x"082082",
   49695 => x"082082",
   49696 => x"082082",
   49697 => x"082082",
   49698 => x"082082",
   49699 => x"082082",
   49700 => x"082082",
   49701 => x"082082",
   49702 => x"082082",
   49703 => x"082082",
   49704 => x"082082",
   49705 => x"082082",
   49706 => x"082082",
   49707 => x"082082",
   49708 => x"082082",
   49709 => x"082082",
   49710 => x"082082",
   49711 => x"082082",
   49712 => x"082082",
   49713 => x"082082",
   49714 => x"082082",
   49715 => x"082041",
   49716 => x"041041",
   49717 => x"041041",
   49718 => x"041041",
   49719 => x"041041",
   49720 => x"041041",
   49721 => x"041041",
   49722 => x"041041",
   49723 => x"041041",
   49724 => x"041041",
   49725 => x"041041",
   49726 => x"041041",
   49727 => x"041041",
   49728 => x"041041",
   49729 => x"041041",
   49730 => x"041041",
   49731 => x"041041",
   49732 => x"041041",
   49733 => x"041041",
   49734 => x"041041",
   49735 => x"041041",
   49736 => x"041041",
   49737 => x"041041",
   49738 => x"041000",
   49739 => x"000000",
   49740 => x"000000",
   49741 => x"000000",
   49742 => x"000000",
   49743 => x"000000",
   49744 => x"000000",
   49745 => x"000000",
   49746 => x"000000",
   49747 => x"000000",
   49748 => x"000000",
   49749 => x"00057f",
   49750 => x"ffffff",
   49751 => x"ffffff",
   49752 => x"ffffff",
   49753 => x"ffffff",
   49754 => x"ffffff",
   49755 => x"ffffff",
   49756 => x"ffffff",
   49757 => x"ffffff",
   49758 => x"ffffff",
   49759 => x"ffffff",
   49760 => x"ffffff",
   49761 => x"ffffff",
   49762 => x"ffffff",
   49763 => x"ffffff",
   49764 => x"ffffff",
   49765 => x"ffffff",
   49766 => x"ffffff",
   49767 => x"ffffff",
   49768 => x"ffffff",
   49769 => x"ffffff",
   49770 => x"ffffff",
   49771 => x"ffffff",
   49772 => x"ffffff",
   49773 => x"ffffff",
   49774 => x"ffffff",
   49775 => x"ffffff",
   49776 => x"ffffff",
   49777 => x"ffffff",
   49778 => x"ffffff",
   49779 => x"ffffff",
   49780 => x"ffffff",
   49781 => x"ffffff",
   49782 => x"ffffff",
   49783 => x"ffffff",
   49784 => x"ffffff",
   49785 => x"ffffff",
   49786 => x"ffffff",
   49787 => x"ffffff",
   49788 => x"ffffff",
   49789 => x"ffffff",
   49790 => x"ffffff",
   49791 => x"ffffff",
   49792 => x"ffffff",
   49793 => x"ffffff",
   49794 => x"ffffff",
   49795 => x"ffffff",
   49796 => x"ffffff",
   49797 => x"ffffff",
   49798 => x"ffffff",
   49799 => x"ffffff",
   49800 => x"ffffff",
   49801 => x"ffffff",
   49802 => x"ffffff",
   49803 => x"ffffff",
   49804 => x"ffffff",
   49805 => x"ffffff",
   49806 => x"ffffff",
   49807 => x"ffffff",
   49808 => x"ffffff",
   49809 => x"ffffff",
   49810 => x"ffffff",
   49811 => x"ffffff",
   49812 => x"ffffff",
   49813 => x"ffffff",
   49814 => x"ffffff",
   49815 => x"ffffff",
   49816 => x"ffffff",
   49817 => x"ffffff",
   49818 => x"ffffff",
   49819 => x"ffffff",
   49820 => x"ffffff",
   49821 => x"ffffff",
   49822 => x"ffffff",
   49823 => x"ffffff",
   49824 => x"ffffff",
   49825 => x"ffffff",
   49826 => x"ffffff",
   49827 => x"ffffff",
   49828 => x"ffffff",
   49829 => x"fffa95",
   49830 => x"abffff",
   49831 => x"ffffff",
   49832 => x"ffffff",
   49833 => x"ffffff",
   49834 => x"ffffff",
   49835 => x"ffffff",
   49836 => x"ffffff",
   49837 => x"ffffff",
   49838 => x"ffffff",
   49839 => x"ffffff",
   49840 => x"ffffff",
   49841 => x"fffac3",
   49842 => x"0c30c3",
   49843 => x"0c30c3",
   49844 => x"0c30c3",
   49845 => x"0c30c3",
   49846 => x"0c30c3",
   49847 => x"0c30c3",
   49848 => x"0c30c3",
   49849 => x"0c30c3",
   49850 => x"0c30c3",
   49851 => x"0c30c3",
   49852 => x"0c30c3",
   49853 => x"082082",
   49854 => x"082082",
   49855 => x"082082",
   49856 => x"082082",
   49857 => x"082082",
   49858 => x"082082",
   49859 => x"082082",
   49860 => x"082082",
   49861 => x"082082",
   49862 => x"082082",
   49863 => x"082082",
   49864 => x"082082",
   49865 => x"082082",
   49866 => x"082082",
   49867 => x"082082",
   49868 => x"082082",
   49869 => x"082082",
   49870 => x"082082",
   49871 => x"082082",
   49872 => x"082082",
   49873 => x"082082",
   49874 => x"082082",
   49875 => x"082041",
   49876 => x"041041",
   49877 => x"041041",
   49878 => x"041041",
   49879 => x"041041",
   49880 => x"041041",
   49881 => x"041041",
   49882 => x"041041",
   49883 => x"041041",
   49884 => x"041041",
   49885 => x"041041",
   49886 => x"041041",
   49887 => x"041041",
   49888 => x"041041",
   49889 => x"041041",
   49890 => x"041041",
   49891 => x"041041",
   49892 => x"041041",
   49893 => x"041041",
   49894 => x"041041",
   49895 => x"041041",
   49896 => x"041041",
   49897 => x"041041",
   49898 => x"041000",
   49899 => x"000000",
   49900 => x"000000",
   49901 => x"000000",
   49902 => x"000000",
   49903 => x"000000",
   49904 => x"000000",
   49905 => x"000000",
   49906 => x"000000",
   49907 => x"000000",
   49908 => x"000000",
   49909 => x"00057f",
   49910 => x"ffffff",
   49911 => x"ffffff",
   49912 => x"ffffff",
   49913 => x"ffffff",
   49914 => x"ffffff",
   49915 => x"ffffff",
   49916 => x"ffffff",
   49917 => x"ffffff",
   49918 => x"ffffff",
   49919 => x"ffffff",
   49920 => x"ffffff",
   49921 => x"ffffff",
   49922 => x"ffffff",
   49923 => x"ffffff",
   49924 => x"ffffff",
   49925 => x"ffffff",
   49926 => x"ffffff",
   49927 => x"ffffff",
   49928 => x"ffffff",
   49929 => x"ffffff",
   49930 => x"ffffff",
   49931 => x"ffffff",
   49932 => x"ffffff",
   49933 => x"ffffff",
   49934 => x"ffffff",
   49935 => x"ffffff",
   49936 => x"ffffff",
   49937 => x"ffffff",
   49938 => x"ffffff",
   49939 => x"ffffff",
   49940 => x"ffffff",
   49941 => x"ffffff",
   49942 => x"ffffff",
   49943 => x"ffffff",
   49944 => x"ffffff",
   49945 => x"ffffff",
   49946 => x"ffffff",
   49947 => x"ffffff",
   49948 => x"ffffff",
   49949 => x"ffffff",
   49950 => x"ffffff",
   49951 => x"ffffff",
   49952 => x"ffffff",
   49953 => x"ffffff",
   49954 => x"ffffff",
   49955 => x"ffffff",
   49956 => x"ffffff",
   49957 => x"ffffff",
   49958 => x"ffffff",
   49959 => x"ffffff",
   49960 => x"ffffff",
   49961 => x"ffffff",
   49962 => x"ffffff",
   49963 => x"ffffff",
   49964 => x"ffffff",
   49965 => x"ffffff",
   49966 => x"ffffff",
   49967 => x"ffffff",
   49968 => x"ffffff",
   49969 => x"ffffff",
   49970 => x"ffffff",
   49971 => x"ffffff",
   49972 => x"ffffff",
   49973 => x"ffffff",
   49974 => x"ffffff",
   49975 => x"ffffff",
   49976 => x"ffffff",
   49977 => x"ffffff",
   49978 => x"ffffff",
   49979 => x"ffffff",
   49980 => x"ffffff",
   49981 => x"ffffff",
   49982 => x"ffffff",
   49983 => x"ffffff",
   49984 => x"ffffff",
   49985 => x"ffffff",
   49986 => x"ffffff",
   49987 => x"ffffff",
   49988 => x"ffffff",
   49989 => x"fffa95",
   49990 => x"abffff",
   49991 => x"ffffff",
   49992 => x"ffffff",
   49993 => x"ffffff",
   49994 => x"ffffff",
   49995 => x"ffffff",
   49996 => x"ffffff",
   49997 => x"ffffff",
   49998 => x"ffffff",
   49999 => x"ffffff",
   50000 => x"ffffff",
   50001 => x"fffac3",
   50002 => x"0c30c3",
   50003 => x"0c30c3",
   50004 => x"0c30c3",
   50005 => x"0c30c3",
   50006 => x"0c30c3",
   50007 => x"0c30c3",
   50008 => x"0c30c3",
   50009 => x"0c30c3",
   50010 => x"0c30c3",
   50011 => x"0c30c3",
   50012 => x"0c30c3",
   50013 => x"082082",
   50014 => x"082082",
   50015 => x"082082",
   50016 => x"082082",
   50017 => x"082082",
   50018 => x"082082",
   50019 => x"082082",
   50020 => x"082082",
   50021 => x"082082",
   50022 => x"082082",
   50023 => x"082082",
   50024 => x"082082",
   50025 => x"082082",
   50026 => x"082082",
   50027 => x"082082",
   50028 => x"082082",
   50029 => x"082082",
   50030 => x"082082",
   50031 => x"082082",
   50032 => x"082082",
   50033 => x"082082",
   50034 => x"082082",
   50035 => x"082041",
   50036 => x"041041",
   50037 => x"041041",
   50038 => x"041041",
   50039 => x"041041",
   50040 => x"041041",
   50041 => x"041041",
   50042 => x"041041",
   50043 => x"041041",
   50044 => x"041041",
   50045 => x"041041",
   50046 => x"041041",
   50047 => x"041041",
   50048 => x"041041",
   50049 => x"041041",
   50050 => x"041041",
   50051 => x"041041",
   50052 => x"041041",
   50053 => x"041041",
   50054 => x"041041",
   50055 => x"041041",
   50056 => x"041041",
   50057 => x"041041",
   50058 => x"041000",
   50059 => x"000000",
   50060 => x"000000",
   50061 => x"000000",
   50062 => x"000000",
   50063 => x"000000",
   50064 => x"000000",
   50065 => x"000000",
   50066 => x"000000",
   50067 => x"000000",
   50068 => x"000000",
   50069 => x"00057f",
   50070 => x"ffffff",
   50071 => x"ffffff",
   50072 => x"ffffff",
   50073 => x"ffffff",
   50074 => x"ffffff",
   50075 => x"ffffff",
   50076 => x"ffffff",
   50077 => x"ffffff",
   50078 => x"ffffff",
   50079 => x"ffffff",
   50080 => x"ffffff",
   50081 => x"ffffff",
   50082 => x"ffffff",
   50083 => x"ffffff",
   50084 => x"ffffff",
   50085 => x"ffffff",
   50086 => x"ffffff",
   50087 => x"ffffff",
   50088 => x"ffffff",
   50089 => x"ffffff",
   50090 => x"ffffff",
   50091 => x"ffffff",
   50092 => x"ffffff",
   50093 => x"ffffff",
   50094 => x"ffffff",
   50095 => x"ffffff",
   50096 => x"ffffff",
   50097 => x"ffffff",
   50098 => x"ffffff",
   50099 => x"ffffff",
   50100 => x"ffffff",
   50101 => x"ffffff",
   50102 => x"ffffff",
   50103 => x"ffffff",
   50104 => x"ffffff",
   50105 => x"ffffff",
   50106 => x"ffffff",
   50107 => x"ffffff",
   50108 => x"ffffff",
   50109 => x"ffffff",
   50110 => x"ffffff",
   50111 => x"ffffff",
   50112 => x"ffffff",
   50113 => x"ffffff",
   50114 => x"ffffff",
   50115 => x"ffffff",
   50116 => x"ffffff",
   50117 => x"ffffff",
   50118 => x"ffffff",
   50119 => x"ffffff",
   50120 => x"ffffff",
   50121 => x"ffffff",
   50122 => x"ffffff",
   50123 => x"ffffff",
   50124 => x"ffffff",
   50125 => x"ffffff",
   50126 => x"ffffff",
   50127 => x"ffffff",
   50128 => x"ffffff",
   50129 => x"ffffff",
   50130 => x"ffffff",
   50131 => x"ffffff",
   50132 => x"ffffff",
   50133 => x"ffffff",
   50134 => x"ffffff",
   50135 => x"ffffff",
   50136 => x"ffffff",
   50137 => x"ffffff",
   50138 => x"ffffff",
   50139 => x"ffffff",
   50140 => x"ffffff",
   50141 => x"ffffff",
   50142 => x"ffffff",
   50143 => x"ffffff",
   50144 => x"ffffff",
   50145 => x"ffffff",
   50146 => x"ffffff",
   50147 => x"ffffff",
   50148 => x"ffffff",
   50149 => x"fffa95",
   50150 => x"abffff",
   50151 => x"ffffff",
   50152 => x"ffffff",
   50153 => x"ffffff",
   50154 => x"ffffff",
   50155 => x"ffffff",
   50156 => x"ffffff",
   50157 => x"ffffff",
   50158 => x"ffffff",
   50159 => x"ffffff",
   50160 => x"ffffff",
   50161 => x"fffac3",
   50162 => x"0c30c3",
   50163 => x"0c30c3",
   50164 => x"0c30c3",
   50165 => x"0c30c3",
   50166 => x"0c30c3",
   50167 => x"0c30c3",
   50168 => x"0c30c3",
   50169 => x"0c30c3",
   50170 => x"0c30c3",
   50171 => x"0c30c3",
   50172 => x"0c30c3",
   50173 => x"082082",
   50174 => x"082082",
   50175 => x"082082",
   50176 => x"082082",
   50177 => x"082082",
   50178 => x"082082",
   50179 => x"082082",
   50180 => x"082082",
   50181 => x"082082",
   50182 => x"082082",
   50183 => x"082082",
   50184 => x"082082",
   50185 => x"082082",
   50186 => x"082082",
   50187 => x"082082",
   50188 => x"082082",
   50189 => x"082082",
   50190 => x"082082",
   50191 => x"082082",
   50192 => x"082082",
   50193 => x"082082",
   50194 => x"082082",
   50195 => x"082041",
   50196 => x"041041",
   50197 => x"041041",
   50198 => x"041041",
   50199 => x"041041",
   50200 => x"041041",
   50201 => x"041041",
   50202 => x"041041",
   50203 => x"041041",
   50204 => x"041041",
   50205 => x"041041",
   50206 => x"041041",
   50207 => x"041041",
   50208 => x"041041",
   50209 => x"041041",
   50210 => x"041041",
   50211 => x"041041",
   50212 => x"041041",
   50213 => x"041041",
   50214 => x"041041",
   50215 => x"041041",
   50216 => x"041041",
   50217 => x"041041",
   50218 => x"041000",
   50219 => x"000000",
   50220 => x"000000",
   50221 => x"000000",
   50222 => x"000000",
   50223 => x"000000",
   50224 => x"000000",
   50225 => x"000000",
   50226 => x"000000",
   50227 => x"000000",
   50228 => x"000000",
   50229 => x"00057f",
   50230 => x"ffffff",
   50231 => x"ffffff",
   50232 => x"ffffff",
   50233 => x"ffffff",
   50234 => x"ffffff",
   50235 => x"ffffff",
   50236 => x"ffffff",
   50237 => x"ffffff",
   50238 => x"ffffff",
   50239 => x"ffffff",
   50240 => x"ffffff",
   50241 => x"ffffff",
   50242 => x"ffffff",
   50243 => x"ffffff",
   50244 => x"ffffff",
   50245 => x"ffffff",
   50246 => x"ffffff",
   50247 => x"ffffff",
   50248 => x"ffffff",
   50249 => x"ffffff",
   50250 => x"ffffff",
   50251 => x"ffffff",
   50252 => x"ffffff",
   50253 => x"ffffff",
   50254 => x"ffffff",
   50255 => x"ffffff",
   50256 => x"ffffff",
   50257 => x"ffffff",
   50258 => x"ffffff",
   50259 => x"ffffff",
   50260 => x"ffffff",
   50261 => x"ffffff",
   50262 => x"ffffff",
   50263 => x"ffffff",
   50264 => x"ffffff",
   50265 => x"ffffff",
   50266 => x"ffffff",
   50267 => x"ffffff",
   50268 => x"ffffff",
   50269 => x"ffffff",
   50270 => x"ffffff",
   50271 => x"ffffff",
   50272 => x"ffffff",
   50273 => x"ffffff",
   50274 => x"ffffff",
   50275 => x"ffffff",
   50276 => x"ffffff",
   50277 => x"ffffff",
   50278 => x"ffffff",
   50279 => x"ffffff",
   50280 => x"ffffff",
   50281 => x"ffffff",
   50282 => x"ffffff",
   50283 => x"ffffff",
   50284 => x"ffffff",
   50285 => x"ffffff",
   50286 => x"ffffff",
   50287 => x"ffffff",
   50288 => x"ffffff",
   50289 => x"ffffff",
   50290 => x"ffffff",
   50291 => x"ffffff",
   50292 => x"ffffff",
   50293 => x"ffffff",
   50294 => x"ffffff",
   50295 => x"ffffff",
   50296 => x"ffffff",
   50297 => x"ffffff",
   50298 => x"ffffff",
   50299 => x"ffffff",
   50300 => x"ffffff",
   50301 => x"ffffff",
   50302 => x"ffffff",
   50303 => x"ffffff",
   50304 => x"ffffff",
   50305 => x"ffffff",
   50306 => x"ffffff",
   50307 => x"ffffff",
   50308 => x"ffffff",
   50309 => x"fffa95",
   50310 => x"abffff",
   50311 => x"ffffff",
   50312 => x"ffffff",
   50313 => x"ffffff",
   50314 => x"ffffff",
   50315 => x"ffffff",
   50316 => x"ffffff",
   50317 => x"ffffff",
   50318 => x"ffffff",
   50319 => x"ffffff",
   50320 => x"ffffff",
   50321 => x"fffac3",
   50322 => x"0c30c3",
   50323 => x"0c30c3",
   50324 => x"0c30c3",
   50325 => x"0c30c3",
   50326 => x"0c30c3",
   50327 => x"0c30c3",
   50328 => x"0c30c3",
   50329 => x"0c30c3",
   50330 => x"0c30c3",
   50331 => x"0c30c3",
   50332 => x"0c30c3",
   50333 => x"082082",
   50334 => x"082082",
   50335 => x"082082",
   50336 => x"082082",
   50337 => x"082082",
   50338 => x"082082",
   50339 => x"082082",
   50340 => x"082082",
   50341 => x"082082",
   50342 => x"082082",
   50343 => x"082082",
   50344 => x"082082",
   50345 => x"082082",
   50346 => x"082082",
   50347 => x"082082",
   50348 => x"082082",
   50349 => x"082082",
   50350 => x"082082",
   50351 => x"082082",
   50352 => x"082082",
   50353 => x"082082",
   50354 => x"082082",
   50355 => x"082041",
   50356 => x"041041",
   50357 => x"041041",
   50358 => x"041041",
   50359 => x"041041",
   50360 => x"041041",
   50361 => x"041041",
   50362 => x"041041",
   50363 => x"041041",
   50364 => x"041041",
   50365 => x"041041",
   50366 => x"041041",
   50367 => x"041041",
   50368 => x"041041",
   50369 => x"041041",
   50370 => x"041041",
   50371 => x"041041",
   50372 => x"041041",
   50373 => x"041041",
   50374 => x"041041",
   50375 => x"041041",
   50376 => x"041041",
   50377 => x"041041",
   50378 => x"041000",
   50379 => x"000000",
   50380 => x"000000",
   50381 => x"000000",
   50382 => x"000000",
   50383 => x"000000",
   50384 => x"000000",
   50385 => x"000000",
   50386 => x"000000",
   50387 => x"000000",
   50388 => x"000000",
   50389 => x"00057f",
   50390 => x"ffffff",
   50391 => x"ffffff",
   50392 => x"ffffff",
   50393 => x"ffffff",
   50394 => x"ffffff",
   50395 => x"ffffff",
   50396 => x"ffffff",
   50397 => x"ffffff",
   50398 => x"ffffff",
   50399 => x"ffffff",
   50400 => x"ffffff",
   50401 => x"ffffff",
   50402 => x"ffffff",
   50403 => x"ffffff",
   50404 => x"ffffff",
   50405 => x"ffffff",
   50406 => x"ffffff",
   50407 => x"ffffff",
   50408 => x"ffffff",
   50409 => x"ffffff",
   50410 => x"ffffff",
   50411 => x"ffffff",
   50412 => x"ffffff",
   50413 => x"ffffff",
   50414 => x"ffffff",
   50415 => x"ffffff",
   50416 => x"ffffff",
   50417 => x"ffffff",
   50418 => x"ffffff",
   50419 => x"ffffff",
   50420 => x"ffffff",
   50421 => x"ffffff",
   50422 => x"ffffff",
   50423 => x"ffffff",
   50424 => x"ffffff",
   50425 => x"ffffff",
   50426 => x"ffffff",
   50427 => x"ffffff",
   50428 => x"ffffff",
   50429 => x"ffffff",
   50430 => x"ffffff",
   50431 => x"ffffff",
   50432 => x"ffffff",
   50433 => x"ffffff",
   50434 => x"ffffff",
   50435 => x"ffffff",
   50436 => x"ffffff",
   50437 => x"ffffff",
   50438 => x"ffffff",
   50439 => x"ffffff",
   50440 => x"ffffff",
   50441 => x"ffffff",
   50442 => x"ffffff",
   50443 => x"ffffff",
   50444 => x"ffffff",
   50445 => x"ffffff",
   50446 => x"ffffff",
   50447 => x"ffffff",
   50448 => x"ffffff",
   50449 => x"ffffff",
   50450 => x"ffffff",
   50451 => x"ffffff",
   50452 => x"ffffff",
   50453 => x"ffffff",
   50454 => x"ffffff",
   50455 => x"ffffff",
   50456 => x"ffffff",
   50457 => x"ffffff",
   50458 => x"ffffff",
   50459 => x"ffffff",
   50460 => x"ffffff",
   50461 => x"ffffff",
   50462 => x"ffffff",
   50463 => x"ffffff",
   50464 => x"ffffff",
   50465 => x"ffffff",
   50466 => x"ffffff",
   50467 => x"ffffff",
   50468 => x"ffffff",
   50469 => x"fffa95",
   50470 => x"abffff",
   50471 => x"ffffff",
   50472 => x"ffffff",
   50473 => x"ffffff",
   50474 => x"ffffff",
   50475 => x"ffffff",
   50476 => x"ffffff",
   50477 => x"ffffff",
   50478 => x"ffffff",
   50479 => x"ffffff",
   50480 => x"ffffff",
   50481 => x"fffac3",
   50482 => x"0c30c3",
   50483 => x"0c30c3",
   50484 => x"0c30c3",
   50485 => x"0c30c3",
   50486 => x"0c30c3",
   50487 => x"0c30c3",
   50488 => x"0c30c3",
   50489 => x"0c30c3",
   50490 => x"0c30c3",
   50491 => x"0c30c3",
   50492 => x"0c30c3",
   50493 => x"082082",
   50494 => x"082082",
   50495 => x"082082",
   50496 => x"082082",
   50497 => x"082082",
   50498 => x"082082",
   50499 => x"082082",
   50500 => x"082082",
   50501 => x"082082",
   50502 => x"082082",
   50503 => x"082082",
   50504 => x"082082",
   50505 => x"082082",
   50506 => x"082082",
   50507 => x"082082",
   50508 => x"082082",
   50509 => x"082082",
   50510 => x"082082",
   50511 => x"082082",
   50512 => x"082082",
   50513 => x"082082",
   50514 => x"082082",
   50515 => x"082041",
   50516 => x"041041",
   50517 => x"041041",
   50518 => x"041041",
   50519 => x"041041",
   50520 => x"041041",
   50521 => x"041041",
   50522 => x"041041",
   50523 => x"041041",
   50524 => x"041041",
   50525 => x"041041",
   50526 => x"041041",
   50527 => x"041041",
   50528 => x"041041",
   50529 => x"041041",
   50530 => x"041041",
   50531 => x"041041",
   50532 => x"041041",
   50533 => x"041041",
   50534 => x"041041",
   50535 => x"041041",
   50536 => x"041041",
   50537 => x"041041",
   50538 => x"041000",
   50539 => x"000000",
   50540 => x"000000",
   50541 => x"000000",
   50542 => x"000000",
   50543 => x"000000",
   50544 => x"000000",
   50545 => x"000000",
   50546 => x"000000",
   50547 => x"000000",
   50548 => x"000000",
   50549 => x"00057f",
   50550 => x"ffffff",
   50551 => x"ffffff",
   50552 => x"ffffff",
   50553 => x"ffffff",
   50554 => x"ffffff",
   50555 => x"ffffff",
   50556 => x"ffffff",
   50557 => x"ffffff",
   50558 => x"ffffff",
   50559 => x"ffffff",
   50560 => x"ffffff",
   50561 => x"ffffff",
   50562 => x"ffffff",
   50563 => x"ffffff",
   50564 => x"ffffff",
   50565 => x"ffffff",
   50566 => x"ffffff",
   50567 => x"ffffff",
   50568 => x"ffffff",
   50569 => x"ffffff",
   50570 => x"ffffff",
   50571 => x"ffffff",
   50572 => x"ffffff",
   50573 => x"ffffff",
   50574 => x"ffffff",
   50575 => x"ffffff",
   50576 => x"ffffff",
   50577 => x"ffffff",
   50578 => x"ffffff",
   50579 => x"ffffff",
   50580 => x"ffffff",
   50581 => x"ffffff",
   50582 => x"ffffff",
   50583 => x"ffffff",
   50584 => x"ffffff",
   50585 => x"ffffff",
   50586 => x"ffffff",
   50587 => x"ffffff",
   50588 => x"ffffff",
   50589 => x"ffffff",
   50590 => x"ffffff",
   50591 => x"ffffff",
   50592 => x"ffffff",
   50593 => x"ffffff",
   50594 => x"ffffff",
   50595 => x"ffffff",
   50596 => x"ffffff",
   50597 => x"ffffff",
   50598 => x"ffffff",
   50599 => x"ffffff",
   50600 => x"ffffff",
   50601 => x"ffffff",
   50602 => x"ffffff",
   50603 => x"ffffff",
   50604 => x"ffffff",
   50605 => x"ffffff",
   50606 => x"ffffff",
   50607 => x"ffffff",
   50608 => x"ffffff",
   50609 => x"ffffff",
   50610 => x"ffffff",
   50611 => x"ffffff",
   50612 => x"ffffff",
   50613 => x"ffffff",
   50614 => x"ffffff",
   50615 => x"ffffff",
   50616 => x"ffffff",
   50617 => x"ffffff",
   50618 => x"ffffff",
   50619 => x"ffffff",
   50620 => x"ffffff",
   50621 => x"ffffff",
   50622 => x"ffffff",
   50623 => x"ffffff",
   50624 => x"ffffff",
   50625 => x"ffffff",
   50626 => x"ffffff",
   50627 => x"ffffff",
   50628 => x"ffffff",
   50629 => x"fffa95",
   50630 => x"abffff",
   50631 => x"ffffff",
   50632 => x"ffffff",
   50633 => x"ffffff",
   50634 => x"ffffff",
   50635 => x"ffffff",
   50636 => x"ffffff",
   50637 => x"ffffff",
   50638 => x"ffffff",
   50639 => x"ffffff",
   50640 => x"ffffff",
   50641 => x"fffac3",
   50642 => x"0c30c3",
   50643 => x"0c30c3",
   50644 => x"0c30c3",
   50645 => x"0c30c3",
   50646 => x"0c30c3",
   50647 => x"0c30c3",
   50648 => x"0c30c3",
   50649 => x"0c30c3",
   50650 => x"0c30c3",
   50651 => x"0c30c3",
   50652 => x"0c30c3",
   50653 => x"082082",
   50654 => x"082082",
   50655 => x"082082",
   50656 => x"082082",
   50657 => x"082082",
   50658 => x"082082",
   50659 => x"082082",
   50660 => x"082082",
   50661 => x"082082",
   50662 => x"082082",
   50663 => x"082082",
   50664 => x"082082",
   50665 => x"082082",
   50666 => x"082082",
   50667 => x"082082",
   50668 => x"082082",
   50669 => x"082082",
   50670 => x"082082",
   50671 => x"082082",
   50672 => x"082082",
   50673 => x"082082",
   50674 => x"082082",
   50675 => x"082041",
   50676 => x"041041",
   50677 => x"041041",
   50678 => x"041041",
   50679 => x"041041",
   50680 => x"041041",
   50681 => x"041041",
   50682 => x"041041",
   50683 => x"041041",
   50684 => x"041041",
   50685 => x"041041",
   50686 => x"041041",
   50687 => x"041041",
   50688 => x"041041",
   50689 => x"041041",
   50690 => x"041041",
   50691 => x"041041",
   50692 => x"041041",
   50693 => x"041041",
   50694 => x"041041",
   50695 => x"041041",
   50696 => x"041041",
   50697 => x"041041",
   50698 => x"041000",
   50699 => x"000000",
   50700 => x"000000",
   50701 => x"000000",
   50702 => x"000000",
   50703 => x"000000",
   50704 => x"000000",
   50705 => x"000000",
   50706 => x"000000",
   50707 => x"000000",
   50708 => x"000000",
   50709 => x"00057f",
   50710 => x"ffffff",
   50711 => x"ffffff",
   50712 => x"ffffff",
   50713 => x"ffffff",
   50714 => x"ffffff",
   50715 => x"ffffff",
   50716 => x"ffffff",
   50717 => x"ffffff",
   50718 => x"ffffff",
   50719 => x"ffffff",
   50720 => x"ffffff",
   50721 => x"ffffff",
   50722 => x"ffffff",
   50723 => x"ffffff",
   50724 => x"ffffff",
   50725 => x"ffffff",
   50726 => x"ffffff",
   50727 => x"ffffff",
   50728 => x"ffffff",
   50729 => x"ffffff",
   50730 => x"ffffff",
   50731 => x"ffffff",
   50732 => x"ffffff",
   50733 => x"ffffff",
   50734 => x"ffffff",
   50735 => x"ffffff",
   50736 => x"ffffff",
   50737 => x"ffffff",
   50738 => x"ffffff",
   50739 => x"ffffff",
   50740 => x"ffffff",
   50741 => x"ffffff",
   50742 => x"ffffff",
   50743 => x"ffffff",
   50744 => x"ffffff",
   50745 => x"ffffff",
   50746 => x"ffffff",
   50747 => x"ffffff",
   50748 => x"ffffff",
   50749 => x"ffffff",
   50750 => x"ffffff",
   50751 => x"ffffff",
   50752 => x"ffffff",
   50753 => x"ffffff",
   50754 => x"ffffff",
   50755 => x"ffffff",
   50756 => x"ffffff",
   50757 => x"ffffff",
   50758 => x"ffffff",
   50759 => x"ffffff",
   50760 => x"ffffff",
   50761 => x"ffffff",
   50762 => x"ffffff",
   50763 => x"ffffff",
   50764 => x"ffffff",
   50765 => x"ffffff",
   50766 => x"ffffff",
   50767 => x"ffffff",
   50768 => x"ffffff",
   50769 => x"ffffff",
   50770 => x"ffffff",
   50771 => x"ffffff",
   50772 => x"ffffff",
   50773 => x"ffffff",
   50774 => x"ffffff",
   50775 => x"ffffff",
   50776 => x"ffffff",
   50777 => x"ffffff",
   50778 => x"ffffff",
   50779 => x"ffffff",
   50780 => x"ffffff",
   50781 => x"ffffff",
   50782 => x"ffffff",
   50783 => x"ffffff",
   50784 => x"ffffff",
   50785 => x"ffffff",
   50786 => x"ffffff",
   50787 => x"ffffff",
   50788 => x"ffffff",
   50789 => x"fffa95",
   50790 => x"abffff",
   50791 => x"ffffff",
   50792 => x"ffffff",
   50793 => x"ffffff",
   50794 => x"ffffff",
   50795 => x"ffffff",
   50796 => x"ffffff",
   50797 => x"ffffff",
   50798 => x"ffffff",
   50799 => x"ffffff",
   50800 => x"ffffff",
   50801 => x"fffac3",
   50802 => x"0c30c3",
   50803 => x"0c30c3",
   50804 => x"0c30c3",
   50805 => x"0c30c3",
   50806 => x"0c30c3",
   50807 => x"0c30c3",
   50808 => x"0c30c3",
   50809 => x"0c30c3",
   50810 => x"0c30c3",
   50811 => x"0c30c3",
   50812 => x"0c30c3",
   50813 => x"082082",
   50814 => x"082082",
   50815 => x"082082",
   50816 => x"082082",
   50817 => x"082082",
   50818 => x"082082",
   50819 => x"082082",
   50820 => x"082082",
   50821 => x"082082",
   50822 => x"082082",
   50823 => x"082082",
   50824 => x"082082",
   50825 => x"082082",
   50826 => x"082082",
   50827 => x"082082",
   50828 => x"082082",
   50829 => x"082082",
   50830 => x"082082",
   50831 => x"082082",
   50832 => x"082082",
   50833 => x"082082",
   50834 => x"082082",
   50835 => x"082041",
   50836 => x"041041",
   50837 => x"041041",
   50838 => x"041041",
   50839 => x"041041",
   50840 => x"041041",
   50841 => x"041041",
   50842 => x"041041",
   50843 => x"041041",
   50844 => x"041041",
   50845 => x"041041",
   50846 => x"041041",
   50847 => x"041041",
   50848 => x"041041",
   50849 => x"041041",
   50850 => x"041041",
   50851 => x"041041",
   50852 => x"041041",
   50853 => x"041041",
   50854 => x"041041",
   50855 => x"041041",
   50856 => x"041041",
   50857 => x"041041",
   50858 => x"041000",
   50859 => x"000000",
   50860 => x"000000",
   50861 => x"000000",
   50862 => x"000000",
   50863 => x"000000",
   50864 => x"000000",
   50865 => x"000000",
   50866 => x"000000",
   50867 => x"000000",
   50868 => x"000000",
   50869 => x"00057f",
   50870 => x"ffffff",
   50871 => x"ffffff",
   50872 => x"ffffff",
   50873 => x"ffffff",
   50874 => x"ffffff",
   50875 => x"ffffff",
   50876 => x"ffffff",
   50877 => x"ffffff",
   50878 => x"ffffff",
   50879 => x"ffffff",
   50880 => x"ffffff",
   50881 => x"ffffff",
   50882 => x"ffffff",
   50883 => x"ffffff",
   50884 => x"ffffff",
   50885 => x"ffffff",
   50886 => x"ffffff",
   50887 => x"ffffff",
   50888 => x"ffffff",
   50889 => x"ffffff",
   50890 => x"ffffff",
   50891 => x"ffffff",
   50892 => x"ffffff",
   50893 => x"ffffff",
   50894 => x"ffffff",
   50895 => x"ffffff",
   50896 => x"ffffff",
   50897 => x"ffffff",
   50898 => x"ffffff",
   50899 => x"ffffff",
   50900 => x"ffffff",
   50901 => x"ffffff",
   50902 => x"ffffff",
   50903 => x"ffffff",
   50904 => x"ffffff",
   50905 => x"ffffff",
   50906 => x"ffffff",
   50907 => x"ffffff",
   50908 => x"ffffff",
   50909 => x"ffffff",
   50910 => x"ffffff",
   50911 => x"ffffff",
   50912 => x"ffffff",
   50913 => x"ffffff",
   50914 => x"ffffff",
   50915 => x"ffffff",
   50916 => x"ffffff",
   50917 => x"ffffff",
   50918 => x"ffffff",
   50919 => x"ffffff",
   50920 => x"ffffff",
   50921 => x"ffffff",
   50922 => x"ffffff",
   50923 => x"ffffff",
   50924 => x"ffffff",
   50925 => x"ffffff",
   50926 => x"ffffff",
   50927 => x"ffffff",
   50928 => x"ffffff",
   50929 => x"ffffff",
   50930 => x"ffffff",
   50931 => x"ffffff",
   50932 => x"ffffff",
   50933 => x"ffffff",
   50934 => x"ffffff",
   50935 => x"ffffff",
   50936 => x"ffffff",
   50937 => x"ffffff",
   50938 => x"ffffff",
   50939 => x"ffffff",
   50940 => x"ffffff",
   50941 => x"ffffff",
   50942 => x"ffffff",
   50943 => x"ffffff",
   50944 => x"ffffff",
   50945 => x"ffffff",
   50946 => x"ffffff",
   50947 => x"ffffff",
   50948 => x"ffffff",
   50949 => x"fffa95",
   50950 => x"abffff",
   50951 => x"ffffff",
   50952 => x"ffffff",
   50953 => x"ffffff",
   50954 => x"ffffff",
   50955 => x"ffffff",
   50956 => x"ffffff",
   50957 => x"ffffff",
   50958 => x"ffffff",
   50959 => x"ffffff",
   50960 => x"ffffff",
   50961 => x"fffac3",
   50962 => x"0c30c3",
   50963 => x"0c30c3",
   50964 => x"0c30c3",
   50965 => x"0c30c3",
   50966 => x"0c30c3",
   50967 => x"0c30c3",
   50968 => x"0c30c3",
   50969 => x"0c30c3",
   50970 => x"0c30c3",
   50971 => x"0c30c3",
   50972 => x"0c30c3",
   50973 => x"082082",
   50974 => x"082082",
   50975 => x"082082",
   50976 => x"082082",
   50977 => x"082082",
   50978 => x"082082",
   50979 => x"082082",
   50980 => x"082082",
   50981 => x"082082",
   50982 => x"082082",
   50983 => x"082082",
   50984 => x"082082",
   50985 => x"082082",
   50986 => x"082082",
   50987 => x"082082",
   50988 => x"082082",
   50989 => x"082082",
   50990 => x"082082",
   50991 => x"082082",
   50992 => x"082082",
   50993 => x"082082",
   50994 => x"082082",
   50995 => x"082041",
   50996 => x"041041",
   50997 => x"041041",
   50998 => x"041041",
   50999 => x"041041",
   51000 => x"041041",
   51001 => x"041041",
   51002 => x"041041",
   51003 => x"041041",
   51004 => x"041041",
   51005 => x"041041",
   51006 => x"041041",
   51007 => x"041041",
   51008 => x"041041",
   51009 => x"041041",
   51010 => x"041041",
   51011 => x"041041",
   51012 => x"041041",
   51013 => x"041041",
   51014 => x"041041",
   51015 => x"041041",
   51016 => x"041041",
   51017 => x"041041",
   51018 => x"041000",
   51019 => x"000000",
   51020 => x"000000",
   51021 => x"000000",
   51022 => x"000000",
   51023 => x"000000",
   51024 => x"000000",
   51025 => x"000000",
   51026 => x"000000",
   51027 => x"000000",
   51028 => x"000000",
   51029 => x"00057f",
   51030 => x"ffffff",
   51031 => x"ffffff",
   51032 => x"ffffff",
   51033 => x"ffffff",
   51034 => x"ffffff",
   51035 => x"ffffff",
   51036 => x"ffffff",
   51037 => x"ffffff",
   51038 => x"ffffff",
   51039 => x"ffffff",
   51040 => x"ffffff",
   51041 => x"ffffff",
   51042 => x"ffffff",
   51043 => x"ffffff",
   51044 => x"ffffff",
   51045 => x"ffffff",
   51046 => x"ffffff",
   51047 => x"ffffff",
   51048 => x"ffffff",
   51049 => x"ffffff",
   51050 => x"ffffff",
   51051 => x"ffffff",
   51052 => x"ffffff",
   51053 => x"ffffff",
   51054 => x"ffffff",
   51055 => x"ffffff",
   51056 => x"ffffff",
   51057 => x"ffffff",
   51058 => x"ffffff",
   51059 => x"ffffff",
   51060 => x"ffffff",
   51061 => x"ffffff",
   51062 => x"ffffff",
   51063 => x"ffffff",
   51064 => x"ffffff",
   51065 => x"ffffff",
   51066 => x"ffffff",
   51067 => x"ffffff",
   51068 => x"ffffff",
   51069 => x"ffffff",
   51070 => x"ffffff",
   51071 => x"ffffff",
   51072 => x"ffffff",
   51073 => x"ffffff",
   51074 => x"ffffff",
   51075 => x"ffffff",
   51076 => x"ffffff",
   51077 => x"ffffff",
   51078 => x"ffffff",
   51079 => x"ffffff",
   51080 => x"ffffff",
   51081 => x"ffffff",
   51082 => x"ffffff",
   51083 => x"ffffff",
   51084 => x"ffffff",
   51085 => x"ffffff",
   51086 => x"ffffff",
   51087 => x"ffffff",
   51088 => x"ffffff",
   51089 => x"ffffff",
   51090 => x"ffffff",
   51091 => x"ffffff",
   51092 => x"ffffff",
   51093 => x"ffffff",
   51094 => x"ffffff",
   51095 => x"ffffff",
   51096 => x"ffffff",
   51097 => x"ffffff",
   51098 => x"ffffff",
   51099 => x"ffffff",
   51100 => x"ffffff",
   51101 => x"ffffff",
   51102 => x"ffffff",
   51103 => x"ffffff",
   51104 => x"ffffff",
   51105 => x"ffffff",
   51106 => x"ffffff",
   51107 => x"ffffff",
   51108 => x"ffffff",
   51109 => x"fffa95",
   51110 => x"abffff",
   51111 => x"ffffff",
   51112 => x"ffffff",
   51113 => x"ffffff",
   51114 => x"ffffff",
   51115 => x"ffffff",
   51116 => x"ffffff",
   51117 => x"ffffff",
   51118 => x"ffffff",
   51119 => x"ffffff",
   51120 => x"ffffff",
   51121 => x"fffac3",
   51122 => x"0c30c3",
   51123 => x"0c30c3",
   51124 => x"0c30c3",
   51125 => x"0c30c3",
   51126 => x"0c30c3",
   51127 => x"0c30c3",
   51128 => x"0c30c3",
   51129 => x"0c30c3",
   51130 => x"0c30c3",
   51131 => x"0c30c3",
   51132 => x"0c30c3",
   51133 => x"082082",
   51134 => x"082082",
   51135 => x"082082",
   51136 => x"082082",
   51137 => x"082082",
   51138 => x"082082",
   51139 => x"082082",
   51140 => x"082082",
   51141 => x"082082",
   51142 => x"082082",
   51143 => x"082082",
   51144 => x"082082",
   51145 => x"082082",
   51146 => x"082082",
   51147 => x"082082",
   51148 => x"082082",
   51149 => x"082082",
   51150 => x"082082",
   51151 => x"082082",
   51152 => x"082082",
   51153 => x"082082",
   51154 => x"082082",
   51155 => x"082041",
   51156 => x"041041",
   51157 => x"041041",
   51158 => x"041041",
   51159 => x"041041",
   51160 => x"041041",
   51161 => x"041041",
   51162 => x"041041",
   51163 => x"041041",
   51164 => x"041041",
   51165 => x"041041",
   51166 => x"041041",
   51167 => x"041041",
   51168 => x"041041",
   51169 => x"041041",
   51170 => x"041041",
   51171 => x"041041",
   51172 => x"041041",
   51173 => x"041041",
   51174 => x"041041",
   51175 => x"041041",
   51176 => x"041041",
   51177 => x"041041",
   51178 => x"041000",
   51179 => x"000000",
   51180 => x"000000",
   51181 => x"000000",
   51182 => x"000000",
   51183 => x"000000",
   51184 => x"000000",
   51185 => x"000000",
   51186 => x"000000",
   51187 => x"000000",
   51188 => x"000000",
   51189 => x"00057f",
   51190 => x"ffffff",
   51191 => x"ffffff",
   51192 => x"ffffff",
   51193 => x"ffffff",
   51194 => x"ffffff",
   51195 => x"ffffff",
   51196 => x"ffffff",
   51197 => x"ffffff",
   51198 => x"ffffff",
   51199 => x"ffffff",
   51200 => x"ffffff",
   51201 => x"ffffff",
   51202 => x"ffffff",
   51203 => x"ffffff",
   51204 => x"ffffff",
   51205 => x"ffffff",
   51206 => x"ffffff",
   51207 => x"ffffff",
   51208 => x"ffffff",
   51209 => x"ffffff",
   51210 => x"ffffff",
   51211 => x"ffffff",
   51212 => x"ffffff",
   51213 => x"ffffff",
   51214 => x"ffffff",
   51215 => x"ffffff",
   51216 => x"ffffff",
   51217 => x"ffffff",
   51218 => x"ffffff",
   51219 => x"ffffff",
   51220 => x"ffffff",
   51221 => x"ffffff",
   51222 => x"ffffff",
   51223 => x"ffffff",
   51224 => x"ffffff",
   51225 => x"ffffff",
   51226 => x"ffffff",
   51227 => x"ffffff",
   51228 => x"ffffff",
   51229 => x"ffffff",
   51230 => x"ffffff",
   51231 => x"ffffff",
   51232 => x"ffffff",
   51233 => x"ffffff",
   51234 => x"ffffff",
   51235 => x"ffffff",
   51236 => x"ffffff",
   51237 => x"ffffff",
   51238 => x"ffffff",
   51239 => x"ffffff",
   51240 => x"ffffff",
   51241 => x"ffffff",
   51242 => x"ffffff",
   51243 => x"ffffff",
   51244 => x"ffffff",
   51245 => x"ffffff",
   51246 => x"ffffff",
   51247 => x"ffffff",
   51248 => x"ffffff",
   51249 => x"ffffff",
   51250 => x"ffffff",
   51251 => x"ffffff",
   51252 => x"ffffff",
   51253 => x"ffffff",
   51254 => x"ffffff",
   51255 => x"ffffff",
   51256 => x"ffffff",
   51257 => x"ffffff",
   51258 => x"ffffff",
   51259 => x"ffffff",
   51260 => x"ffffff",
   51261 => x"ffffff",
   51262 => x"ffffff",
   51263 => x"ffffff",
   51264 => x"ffffff",
   51265 => x"ffffff",
   51266 => x"ffffff",
   51267 => x"ffffff",
   51268 => x"ffffff",
   51269 => x"fffa95",
   51270 => x"abffff",
   51271 => x"ffffff",
   51272 => x"ffffff",
   51273 => x"ffffff",
   51274 => x"ffffff",
   51275 => x"ffffff",
   51276 => x"ffffff",
   51277 => x"ffffff",
   51278 => x"ffffff",
   51279 => x"ffffff",
   51280 => x"ffffff",
   51281 => x"fffac3",
   51282 => x"0c30c3",
   51283 => x"0c30c3",
   51284 => x"0c30c3",
   51285 => x"0c30c3",
   51286 => x"0c30c3",
   51287 => x"0c30c3",
   51288 => x"0c30c3",
   51289 => x"0c30c3",
   51290 => x"0c30c3",
   51291 => x"0c30c3",
   51292 => x"0c30c3",
   51293 => x"082082",
   51294 => x"082082",
   51295 => x"082082",
   51296 => x"082082",
   51297 => x"082082",
   51298 => x"082082",
   51299 => x"082082",
   51300 => x"082082",
   51301 => x"082082",
   51302 => x"082082",
   51303 => x"082082",
   51304 => x"082082",
   51305 => x"082082",
   51306 => x"082082",
   51307 => x"082082",
   51308 => x"082082",
   51309 => x"082082",
   51310 => x"082082",
   51311 => x"082082",
   51312 => x"082082",
   51313 => x"082082",
   51314 => x"082082",
   51315 => x"082041",
   51316 => x"041041",
   51317 => x"041041",
   51318 => x"041041",
   51319 => x"041041",
   51320 => x"041041",
   51321 => x"041041",
   51322 => x"041041",
   51323 => x"041041",
   51324 => x"041041",
   51325 => x"041041",
   51326 => x"041041",
   51327 => x"041041",
   51328 => x"041041",
   51329 => x"041041",
   51330 => x"041041",
   51331 => x"041041",
   51332 => x"041041",
   51333 => x"041041",
   51334 => x"041041",
   51335 => x"041041",
   51336 => x"041041",
   51337 => x"041041",
   51338 => x"041000",
   51339 => x"000000",
   51340 => x"000000",
   51341 => x"000000",
   51342 => x"000000",
   51343 => x"000000",
   51344 => x"000000",
   51345 => x"000000",
   51346 => x"000000",
   51347 => x"000000",
   51348 => x"000000",
   51349 => x"00057f",
   51350 => x"ffffff",
   51351 => x"ffffff",
   51352 => x"ffffff",
   51353 => x"ffffea",
   51354 => x"aaaaaa",
   51355 => x"aaaaaa",
   51356 => x"aaaaaa",
   51357 => x"ffffff",
   51358 => x"ffffff",
   51359 => x"ffffff",
   51360 => x"ffffff",
   51361 => x"ffffff",
   51362 => x"ffffff",
   51363 => x"ffffff",
   51364 => x"ffffff",
   51365 => x"ffffff",
   51366 => x"ffffff",
   51367 => x"ffffff",
   51368 => x"ffffff",
   51369 => x"ffffff",
   51370 => x"ffffff",
   51371 => x"ffffff",
   51372 => x"ffffff",
   51373 => x"ffffff",
   51374 => x"ffffff",
   51375 => x"ffffff",
   51376 => x"ffffff",
   51377 => x"ffffff",
   51378 => x"ffffff",
   51379 => x"ffffff",
   51380 => x"ffffff",
   51381 => x"ffffff",
   51382 => x"ffffff",
   51383 => x"ffffff",
   51384 => x"ffffff",
   51385 => x"ffffff",
   51386 => x"ffffff",
   51387 => x"ffffff",
   51388 => x"ffffff",
   51389 => x"ffffff",
   51390 => x"ffffff",
   51391 => x"ffffff",
   51392 => x"ffffff",
   51393 => x"ffffff",
   51394 => x"ffffff",
   51395 => x"ffffff",
   51396 => x"ffffff",
   51397 => x"ffffff",
   51398 => x"ffffff",
   51399 => x"ffffff",
   51400 => x"ffffff",
   51401 => x"ffffff",
   51402 => x"ffffff",
   51403 => x"ffffff",
   51404 => x"ffffff",
   51405 => x"ffffff",
   51406 => x"ffffff",
   51407 => x"ffffff",
   51408 => x"ffffff",
   51409 => x"ffffff",
   51410 => x"ffffff",
   51411 => x"ffffff",
   51412 => x"ffffff",
   51413 => x"ffffff",
   51414 => x"ffffff",
   51415 => x"ffffff",
   51416 => x"ffffff",
   51417 => x"ffffff",
   51418 => x"ffffff",
   51419 => x"ffffff",
   51420 => x"ffffff",
   51421 => x"ffffff",
   51422 => x"ffffff",
   51423 => x"ffffff",
   51424 => x"ffffff",
   51425 => x"ffffff",
   51426 => x"ffffff",
   51427 => x"ffffff",
   51428 => x"ffffff",
   51429 => x"fffa95",
   51430 => x"abffff",
   51431 => x"ffffff",
   51432 => x"ffffff",
   51433 => x"ffffff",
   51434 => x"ffffff",
   51435 => x"ffffff",
   51436 => x"ffffff",
   51437 => x"ffffff",
   51438 => x"ffffff",
   51439 => x"ffffff",
   51440 => x"ffffff",
   51441 => x"fffac3",
   51442 => x"0c30c3",
   51443 => x"0c30c3",
   51444 => x"0c30c3",
   51445 => x"0c30c3",
   51446 => x"0c30c3",
   51447 => x"0c30c3",
   51448 => x"0c30c3",
   51449 => x"0c30c3",
   51450 => x"0c30c3",
   51451 => x"0c30c3",
   51452 => x"0c30c3",
   51453 => x"082082",
   51454 => x"082082",
   51455 => x"082082",
   51456 => x"082082",
   51457 => x"082082",
   51458 => x"082082",
   51459 => x"082082",
   51460 => x"082082",
   51461 => x"082082",
   51462 => x"082082",
   51463 => x"082082",
   51464 => x"082082",
   51465 => x"082082",
   51466 => x"082082",
   51467 => x"082082",
   51468 => x"082082",
   51469 => x"082082",
   51470 => x"082082",
   51471 => x"082082",
   51472 => x"082082",
   51473 => x"082082",
   51474 => x"082082",
   51475 => x"082041",
   51476 => x"041041",
   51477 => x"041041",
   51478 => x"041041",
   51479 => x"041041",
   51480 => x"041041",
   51481 => x"041041",
   51482 => x"041041",
   51483 => x"041041",
   51484 => x"041041",
   51485 => x"041041",
   51486 => x"041041",
   51487 => x"041041",
   51488 => x"041041",
   51489 => x"041041",
   51490 => x"041041",
   51491 => x"041041",
   51492 => x"041041",
   51493 => x"041041",
   51494 => x"041041",
   51495 => x"041041",
   51496 => x"041041",
   51497 => x"041041",
   51498 => x"041000",
   51499 => x"000000",
   51500 => x"000000",
   51501 => x"000000",
   51502 => x"000000",
   51503 => x"000000",
   51504 => x"000000",
   51505 => x"000000",
   51506 => x"000000",
   51507 => x"000000",
   51508 => x"000000",
   51509 => x"00057f",
   51510 => x"ffffff",
   51511 => x"ffffff",
   51512 => x"ffffff",
   51513 => x"ffffd5",
   51514 => x"000000",
   51515 => x"000000",
   51516 => x"000000",
   51517 => x"55556a",
   51518 => x"ffffff",
   51519 => x"ffffff",
   51520 => x"ffffff",
   51521 => x"ffffff",
   51522 => x"ffffff",
   51523 => x"ffffff",
   51524 => x"ffffff",
   51525 => x"ffffff",
   51526 => x"ffffff",
   51527 => x"ffffff",
   51528 => x"ffffff",
   51529 => x"ffffff",
   51530 => x"ffffff",
   51531 => x"ffffff",
   51532 => x"ffffff",
   51533 => x"ffffff",
   51534 => x"ffffff",
   51535 => x"ffffff",
   51536 => x"ffffff",
   51537 => x"ffffff",
   51538 => x"ffffff",
   51539 => x"ffffff",
   51540 => x"ffffff",
   51541 => x"ffffff",
   51542 => x"ffffff",
   51543 => x"ffffff",
   51544 => x"ffffff",
   51545 => x"ffffff",
   51546 => x"ffffff",
   51547 => x"ffffff",
   51548 => x"ffffff",
   51549 => x"ffffff",
   51550 => x"ffffff",
   51551 => x"ffffff",
   51552 => x"ffffff",
   51553 => x"ffffff",
   51554 => x"ffffff",
   51555 => x"ffffff",
   51556 => x"ffffff",
   51557 => x"ffffff",
   51558 => x"ffffff",
   51559 => x"ffffff",
   51560 => x"ffffff",
   51561 => x"ffffff",
   51562 => x"ffffff",
   51563 => x"ffffff",
   51564 => x"ffffff",
   51565 => x"ffffff",
   51566 => x"ffffff",
   51567 => x"ffffff",
   51568 => x"ffffff",
   51569 => x"ffffff",
   51570 => x"ffffff",
   51571 => x"ffffff",
   51572 => x"ffffff",
   51573 => x"ffffff",
   51574 => x"ffffff",
   51575 => x"ffffff",
   51576 => x"ffffff",
   51577 => x"ffffff",
   51578 => x"ffffff",
   51579 => x"ffffff",
   51580 => x"ffffff",
   51581 => x"ffffff",
   51582 => x"ffffff",
   51583 => x"ffffff",
   51584 => x"ffffff",
   51585 => x"ffffff",
   51586 => x"ffffff",
   51587 => x"ffffff",
   51588 => x"ffffff",
   51589 => x"fffa95",
   51590 => x"abffff",
   51591 => x"ffffff",
   51592 => x"ffffff",
   51593 => x"ffffff",
   51594 => x"ffffff",
   51595 => x"ffffff",
   51596 => x"ffffff",
   51597 => x"ffffff",
   51598 => x"ffffff",
   51599 => x"ffffff",
   51600 => x"ffffff",
   51601 => x"fffac3",
   51602 => x"0c30c3",
   51603 => x"0c30c3",
   51604 => x"0c30c3",
   51605 => x"0c30c3",
   51606 => x"0c30c3",
   51607 => x"0c30c3",
   51608 => x"0c30c3",
   51609 => x"0c30c3",
   51610 => x"0c30c3",
   51611 => x"0c30c3",
   51612 => x"0c30c3",
   51613 => x"082082",
   51614 => x"082082",
   51615 => x"082082",
   51616 => x"082082",
   51617 => x"082082",
   51618 => x"082082",
   51619 => x"082082",
   51620 => x"082082",
   51621 => x"082082",
   51622 => x"082082",
   51623 => x"082082",
   51624 => x"082082",
   51625 => x"082082",
   51626 => x"082082",
   51627 => x"082082",
   51628 => x"082082",
   51629 => x"082082",
   51630 => x"082082",
   51631 => x"082082",
   51632 => x"082082",
   51633 => x"082082",
   51634 => x"082082",
   51635 => x"082041",
   51636 => x"041041",
   51637 => x"041041",
   51638 => x"041041",
   51639 => x"041041",
   51640 => x"041041",
   51641 => x"041041",
   51642 => x"041041",
   51643 => x"041041",
   51644 => x"041041",
   51645 => x"041041",
   51646 => x"041041",
   51647 => x"041041",
   51648 => x"041041",
   51649 => x"041041",
   51650 => x"041041",
   51651 => x"041041",
   51652 => x"041041",
   51653 => x"041041",
   51654 => x"041041",
   51655 => x"041041",
   51656 => x"041041",
   51657 => x"041041",
   51658 => x"041000",
   51659 => x"000000",
   51660 => x"000000",
   51661 => x"000000",
   51662 => x"000000",
   51663 => x"000000",
   51664 => x"000000",
   51665 => x"000000",
   51666 => x"000000",
   51667 => x"000000",
   51668 => x"000000",
   51669 => x"00057f",
   51670 => x"ffffff",
   51671 => x"ffffff",
   51672 => x"ffffff",
   51673 => x"ffffd5",
   51674 => x"000000",
   51675 => x"000000",
   51676 => x"000000",
   51677 => x"000000",
   51678 => x"57ffff",
   51679 => x"ffffff",
   51680 => x"ffffff",
   51681 => x"ffffff",
   51682 => x"ffffff",
   51683 => x"ffffff",
   51684 => x"ffffff",
   51685 => x"ffffff",
   51686 => x"ffffff",
   51687 => x"ffffff",
   51688 => x"ffffff",
   51689 => x"ffffff",
   51690 => x"ffffff",
   51691 => x"ffffff",
   51692 => x"ffffff",
   51693 => x"ffffff",
   51694 => x"ffffff",
   51695 => x"ffffff",
   51696 => x"ffffff",
   51697 => x"ffffff",
   51698 => x"ffffff",
   51699 => x"ffffff",
   51700 => x"ffffff",
   51701 => x"ffffff",
   51702 => x"ffffff",
   51703 => x"ffffff",
   51704 => x"ffffff",
   51705 => x"ffffff",
   51706 => x"ffffff",
   51707 => x"ffffff",
   51708 => x"ffffff",
   51709 => x"ffffff",
   51710 => x"ffffff",
   51711 => x"ffffff",
   51712 => x"ffffff",
   51713 => x"ffffff",
   51714 => x"ffffff",
   51715 => x"ffffff",
   51716 => x"ffffff",
   51717 => x"ffffff",
   51718 => x"ffffff",
   51719 => x"ffffff",
   51720 => x"ffffff",
   51721 => x"ffffff",
   51722 => x"ffffff",
   51723 => x"ffffff",
   51724 => x"ffffff",
   51725 => x"ffffff",
   51726 => x"ffffff",
   51727 => x"ffffff",
   51728 => x"ffffff",
   51729 => x"ffffff",
   51730 => x"ffffff",
   51731 => x"ffffff",
   51732 => x"ffffff",
   51733 => x"ffffff",
   51734 => x"ffffff",
   51735 => x"ffffff",
   51736 => x"ffffff",
   51737 => x"ffffff",
   51738 => x"ffffff",
   51739 => x"ffffff",
   51740 => x"ffffff",
   51741 => x"ffffff",
   51742 => x"ffffff",
   51743 => x"ffffff",
   51744 => x"ffffff",
   51745 => x"ffffff",
   51746 => x"ffffff",
   51747 => x"ffffff",
   51748 => x"ffffff",
   51749 => x"fffa95",
   51750 => x"abffff",
   51751 => x"ffffff",
   51752 => x"ffffff",
   51753 => x"ffffff",
   51754 => x"ffffff",
   51755 => x"ffffff",
   51756 => x"ffffff",
   51757 => x"ffffff",
   51758 => x"ffffff",
   51759 => x"ffffff",
   51760 => x"ffffff",
   51761 => x"fffac3",
   51762 => x"0c30c3",
   51763 => x"0c30c3",
   51764 => x"0c30c3",
   51765 => x"0c30c3",
   51766 => x"0c30c3",
   51767 => x"0c30c3",
   51768 => x"0c30c3",
   51769 => x"0c30c3",
   51770 => x"0c30c3",
   51771 => x"0c30c3",
   51772 => x"0c30c3",
   51773 => x"082082",
   51774 => x"082082",
   51775 => x"082082",
   51776 => x"082082",
   51777 => x"082082",
   51778 => x"082082",
   51779 => x"082082",
   51780 => x"082082",
   51781 => x"082082",
   51782 => x"082082",
   51783 => x"082082",
   51784 => x"082082",
   51785 => x"082082",
   51786 => x"082082",
   51787 => x"082082",
   51788 => x"082082",
   51789 => x"082082",
   51790 => x"082082",
   51791 => x"082082",
   51792 => x"082082",
   51793 => x"082082",
   51794 => x"082082",
   51795 => x"082041",
   51796 => x"041041",
   51797 => x"041041",
   51798 => x"041041",
   51799 => x"041041",
   51800 => x"041041",
   51801 => x"041041",
   51802 => x"041041",
   51803 => x"041041",
   51804 => x"041041",
   51805 => x"041041",
   51806 => x"041041",
   51807 => x"041041",
   51808 => x"041041",
   51809 => x"041041",
   51810 => x"041041",
   51811 => x"041041",
   51812 => x"041041",
   51813 => x"041041",
   51814 => x"041041",
   51815 => x"041041",
   51816 => x"041041",
   51817 => x"041041",
   51818 => x"041000",
   51819 => x"000000",
   51820 => x"000000",
   51821 => x"000000",
   51822 => x"000000",
   51823 => x"000000",
   51824 => x"000000",
   51825 => x"000000",
   51826 => x"000000",
   51827 => x"000000",
   51828 => x"000000",
   51829 => x"00057f",
   51830 => x"ffffff",
   51831 => x"ffffff",
   51832 => x"ffffff",
   51833 => x"ffffd5",
   51834 => x"000000",
   51835 => x"000000",
   51836 => x"000000",
   51837 => x"000000",
   51838 => x"015fff",
   51839 => x"ffffff",
   51840 => x"ffffff",
   51841 => x"ffffff",
   51842 => x"ffffff",
   51843 => x"ffffff",
   51844 => x"ffffff",
   51845 => x"ffffff",
   51846 => x"ffffff",
   51847 => x"ffffff",
   51848 => x"ffffff",
   51849 => x"ffffff",
   51850 => x"ffffff",
   51851 => x"ffffff",
   51852 => x"ffffff",
   51853 => x"ffffff",
   51854 => x"ffffff",
   51855 => x"ffffff",
   51856 => x"ffffff",
   51857 => x"ffffff",
   51858 => x"ffffff",
   51859 => x"ffffff",
   51860 => x"ffffff",
   51861 => x"ffffff",
   51862 => x"ffffff",
   51863 => x"ffffff",
   51864 => x"ffffff",
   51865 => x"ffffff",
   51866 => x"ffffff",
   51867 => x"ffffff",
   51868 => x"ffffff",
   51869 => x"ffffff",
   51870 => x"ffffff",
   51871 => x"ffffff",
   51872 => x"ffffff",
   51873 => x"ffffff",
   51874 => x"ffffff",
   51875 => x"ffffff",
   51876 => x"ffffff",
   51877 => x"ffffff",
   51878 => x"ffffff",
   51879 => x"ffffff",
   51880 => x"ffffff",
   51881 => x"ffffff",
   51882 => x"ffffff",
   51883 => x"ffffff",
   51884 => x"ffffff",
   51885 => x"ffffff",
   51886 => x"ffffff",
   51887 => x"ffffff",
   51888 => x"ffffff",
   51889 => x"ffffff",
   51890 => x"ffffff",
   51891 => x"ffffff",
   51892 => x"ffffff",
   51893 => x"ffffff",
   51894 => x"ffffff",
   51895 => x"ffffff",
   51896 => x"ffffff",
   51897 => x"ffffff",
   51898 => x"ffffff",
   51899 => x"ffffff",
   51900 => x"ffffff",
   51901 => x"ffffff",
   51902 => x"ffffff",
   51903 => x"ffffff",
   51904 => x"ffffff",
   51905 => x"ffffff",
   51906 => x"ffffff",
   51907 => x"ffffff",
   51908 => x"ffffff",
   51909 => x"fffa95",
   51910 => x"abffff",
   51911 => x"ffffff",
   51912 => x"ffffff",
   51913 => x"ffffff",
   51914 => x"ffffff",
   51915 => x"ffffff",
   51916 => x"ffffff",
   51917 => x"ffffff",
   51918 => x"ffffff",
   51919 => x"ffffff",
   51920 => x"ffffff",
   51921 => x"fffac3",
   51922 => x"0c30c3",
   51923 => x"0c30c3",
   51924 => x"0c30c3",
   51925 => x"0c30c3",
   51926 => x"0c30c3",
   51927 => x"0c30c3",
   51928 => x"0c30c3",
   51929 => x"0c30c3",
   51930 => x"0c30c3",
   51931 => x"0c30c3",
   51932 => x"0c30c3",
   51933 => x"082082",
   51934 => x"082082",
   51935 => x"082082",
   51936 => x"082082",
   51937 => x"082082",
   51938 => x"082082",
   51939 => x"082082",
   51940 => x"082082",
   51941 => x"082082",
   51942 => x"082082",
   51943 => x"082082",
   51944 => x"082082",
   51945 => x"082082",
   51946 => x"082082",
   51947 => x"082082",
   51948 => x"082082",
   51949 => x"082082",
   51950 => x"082082",
   51951 => x"082082",
   51952 => x"082082",
   51953 => x"082082",
   51954 => x"082082",
   51955 => x"082041",
   51956 => x"041041",
   51957 => x"041041",
   51958 => x"041041",
   51959 => x"041041",
   51960 => x"041041",
   51961 => x"041041",
   51962 => x"041041",
   51963 => x"041041",
   51964 => x"041041",
   51965 => x"041041",
   51966 => x"041041",
   51967 => x"041041",
   51968 => x"041041",
   51969 => x"041041",
   51970 => x"041041",
   51971 => x"041041",
   51972 => x"041041",
   51973 => x"041041",
   51974 => x"041041",
   51975 => x"041041",
   51976 => x"041041",
   51977 => x"041041",
   51978 => x"041000",
   51979 => x"000000",
   51980 => x"000000",
   51981 => x"000000",
   51982 => x"000000",
   51983 => x"000000",
   51984 => x"000000",
   51985 => x"000000",
   51986 => x"000000",
   51987 => x"000000",
   51988 => x"000000",
   51989 => x"00057f",
   51990 => x"ffffff",
   51991 => x"ffffff",
   51992 => x"ffffff",
   51993 => x"ffffd5",
   51994 => x"000015",
   51995 => x"aaaaaa",
   51996 => x"aaaaaa",
   51997 => x"555000",
   51998 => x"00057f",
   51999 => x"ffffff",
   52000 => x"ffffff",
   52001 => x"ffffff",
   52002 => x"ffffff",
   52003 => x"ffffff",
   52004 => x"ffffff",
   52005 => x"ffffff",
   52006 => x"ffffff",
   52007 => x"ffffff",
   52008 => x"ffffff",
   52009 => x"ffffff",
   52010 => x"ffffff",
   52011 => x"ffffff",
   52012 => x"ffffff",
   52013 => x"ffffff",
   52014 => x"ffffff",
   52015 => x"ffffff",
   52016 => x"ffffff",
   52017 => x"ffffff",
   52018 => x"ffffff",
   52019 => x"ffffff",
   52020 => x"ffffff",
   52021 => x"ffffff",
   52022 => x"ffffff",
   52023 => x"ffffff",
   52024 => x"ffffff",
   52025 => x"ffffff",
   52026 => x"ffffff",
   52027 => x"ffffff",
   52028 => x"ffffff",
   52029 => x"ffffff",
   52030 => x"ffffff",
   52031 => x"ffffff",
   52032 => x"ffffff",
   52033 => x"ffffff",
   52034 => x"ffffff",
   52035 => x"ffffff",
   52036 => x"ffffff",
   52037 => x"ffffff",
   52038 => x"ffffff",
   52039 => x"ffffff",
   52040 => x"ffffff",
   52041 => x"ffffff",
   52042 => x"ffffff",
   52043 => x"ffffff",
   52044 => x"ffffff",
   52045 => x"ffffff",
   52046 => x"ffffff",
   52047 => x"ffffff",
   52048 => x"ffffff",
   52049 => x"ffffff",
   52050 => x"ffffff",
   52051 => x"ffffff",
   52052 => x"ffffff",
   52053 => x"ffffff",
   52054 => x"ffffff",
   52055 => x"ffffff",
   52056 => x"ffffff",
   52057 => x"ffffff",
   52058 => x"ffffff",
   52059 => x"ffffff",
   52060 => x"ffffff",
   52061 => x"ffffff",
   52062 => x"ffffff",
   52063 => x"ffffff",
   52064 => x"ffffff",
   52065 => x"ffffff",
   52066 => x"ffffff",
   52067 => x"ffffff",
   52068 => x"ffffff",
   52069 => x"fffa95",
   52070 => x"abffff",
   52071 => x"ffffff",
   52072 => x"ffffff",
   52073 => x"ffffff",
   52074 => x"ffffff",
   52075 => x"ffffff",
   52076 => x"ffffff",
   52077 => x"ffffff",
   52078 => x"ffffff",
   52079 => x"ffffff",
   52080 => x"ffffff",
   52081 => x"fffac3",
   52082 => x"0c30c3",
   52083 => x"0c30c3",
   52084 => x"0c30c3",
   52085 => x"0c30c3",
   52086 => x"0c30c3",
   52087 => x"0c30c3",
   52088 => x"0c30c3",
   52089 => x"0c30c3",
   52090 => x"0c30c3",
   52091 => x"0c30c3",
   52092 => x"0c30c3",
   52093 => x"082082",
   52094 => x"082082",
   52095 => x"082082",
   52096 => x"082082",
   52097 => x"082082",
   52098 => x"082082",
   52099 => x"082082",
   52100 => x"082082",
   52101 => x"082082",
   52102 => x"082082",
   52103 => x"082082",
   52104 => x"082082",
   52105 => x"082082",
   52106 => x"082082",
   52107 => x"082082",
   52108 => x"082082",
   52109 => x"082082",
   52110 => x"082082",
   52111 => x"082082",
   52112 => x"082082",
   52113 => x"082082",
   52114 => x"082082",
   52115 => x"082041",
   52116 => x"041041",
   52117 => x"041041",
   52118 => x"041041",
   52119 => x"041041",
   52120 => x"041041",
   52121 => x"041041",
   52122 => x"041041",
   52123 => x"041041",
   52124 => x"041041",
   52125 => x"041041",
   52126 => x"041041",
   52127 => x"041041",
   52128 => x"041041",
   52129 => x"041041",
   52130 => x"041041",
   52131 => x"041041",
   52132 => x"041041",
   52133 => x"041041",
   52134 => x"041041",
   52135 => x"041041",
   52136 => x"041041",
   52137 => x"041041",
   52138 => x"041000",
   52139 => x"000000",
   52140 => x"000000",
   52141 => x"000000",
   52142 => x"000000",
   52143 => x"000000",
   52144 => x"000000",
   52145 => x"000000",
   52146 => x"000000",
   52147 => x"000000",
   52148 => x"000000",
   52149 => x"00057f",
   52150 => x"ffffff",
   52151 => x"ffffff",
   52152 => x"ffffff",
   52153 => x"ffffd5",
   52154 => x"00002a",
   52155 => x"ffffff",
   52156 => x"ffffff",
   52157 => x"fea540",
   52158 => x"00057f",
   52159 => x"ffffff",
   52160 => x"ffffff",
   52161 => x"ffffff",
   52162 => x"ffffff",
   52163 => x"ffffff",
   52164 => x"ffffff",
   52165 => x"ffffff",
   52166 => x"ffffff",
   52167 => x"ffffff",
   52168 => x"ffffff",
   52169 => x"ffffff",
   52170 => x"ffffff",
   52171 => x"ffffff",
   52172 => x"ffffff",
   52173 => x"ffffff",
   52174 => x"ffffff",
   52175 => x"ffffff",
   52176 => x"ffffff",
   52177 => x"ffffff",
   52178 => x"ffffff",
   52179 => x"ffffff",
   52180 => x"ffffff",
   52181 => x"ffffff",
   52182 => x"ffffff",
   52183 => x"ffffff",
   52184 => x"ffffff",
   52185 => x"ffffff",
   52186 => x"ffffff",
   52187 => x"ffffff",
   52188 => x"ffffff",
   52189 => x"ffffff",
   52190 => x"ffffff",
   52191 => x"ffffff",
   52192 => x"ffffff",
   52193 => x"ffffff",
   52194 => x"ffffff",
   52195 => x"ffffff",
   52196 => x"ffffff",
   52197 => x"ffffff",
   52198 => x"ffffff",
   52199 => x"ffffff",
   52200 => x"ffffff",
   52201 => x"ffffff",
   52202 => x"ffffff",
   52203 => x"ffffff",
   52204 => x"ffffff",
   52205 => x"ffffff",
   52206 => x"ffffff",
   52207 => x"ffffff",
   52208 => x"ffffff",
   52209 => x"ffffff",
   52210 => x"ffffff",
   52211 => x"ffffff",
   52212 => x"ffffff",
   52213 => x"ffffff",
   52214 => x"ffffff",
   52215 => x"ffffff",
   52216 => x"ffffff",
   52217 => x"ffffff",
   52218 => x"ffffff",
   52219 => x"ffffff",
   52220 => x"ffffff",
   52221 => x"ffffff",
   52222 => x"ffffff",
   52223 => x"ffffff",
   52224 => x"ffffff",
   52225 => x"ffffff",
   52226 => x"ffffff",
   52227 => x"ffffff",
   52228 => x"ffffff",
   52229 => x"fffa95",
   52230 => x"abffff",
   52231 => x"ffffff",
   52232 => x"ffffff",
   52233 => x"ffffff",
   52234 => x"ffffff",
   52235 => x"ffffff",
   52236 => x"ffffff",
   52237 => x"ffffff",
   52238 => x"ffffff",
   52239 => x"ffffff",
   52240 => x"ffffff",
   52241 => x"fffac3",
   52242 => x"0c30c3",
   52243 => x"0c30c3",
   52244 => x"0c30c3",
   52245 => x"0c30c3",
   52246 => x"0c30c3",
   52247 => x"0c30c3",
   52248 => x"0c30c3",
   52249 => x"0c30c3",
   52250 => x"0c30c3",
   52251 => x"0c30c3",
   52252 => x"0c30c3",
   52253 => x"082082",
   52254 => x"082082",
   52255 => x"082082",
   52256 => x"082082",
   52257 => x"082082",
   52258 => x"082082",
   52259 => x"082082",
   52260 => x"082082",
   52261 => x"082082",
   52262 => x"082082",
   52263 => x"082082",
   52264 => x"082082",
   52265 => x"082082",
   52266 => x"082082",
   52267 => x"082082",
   52268 => x"082082",
   52269 => x"082082",
   52270 => x"082082",
   52271 => x"082082",
   52272 => x"082082",
   52273 => x"082082",
   52274 => x"082082",
   52275 => x"082041",
   52276 => x"041041",
   52277 => x"041041",
   52278 => x"041041",
   52279 => x"041041",
   52280 => x"041041",
   52281 => x"041041",
   52282 => x"041041",
   52283 => x"041041",
   52284 => x"041041",
   52285 => x"041041",
   52286 => x"041041",
   52287 => x"041041",
   52288 => x"041041",
   52289 => x"041041",
   52290 => x"041041",
   52291 => x"041041",
   52292 => x"041041",
   52293 => x"041041",
   52294 => x"041041",
   52295 => x"041041",
   52296 => x"041041",
   52297 => x"041041",
   52298 => x"041000",
   52299 => x"000000",
   52300 => x"000000",
   52301 => x"000000",
   52302 => x"000000",
   52303 => x"000000",
   52304 => x"000000",
   52305 => x"000000",
   52306 => x"000000",
   52307 => x"000000",
   52308 => x"000000",
   52309 => x"00057f",
   52310 => x"ffffff",
   52311 => x"ffffff",
   52312 => x"ffffff",
   52313 => x"ffffd5",
   52314 => x"00002a",
   52315 => x"ffffff",
   52316 => x"ffffff",
   52317 => x"fffa80",
   52318 => x"00002a",
   52319 => x"ffffff",
   52320 => x"ffffff",
   52321 => x"ffffff",
   52322 => x"ffffff",
   52323 => x"ffffff",
   52324 => x"ffffff",
   52325 => x"ffffff",
   52326 => x"ffffff",
   52327 => x"ffffff",
   52328 => x"ffffff",
   52329 => x"ffffff",
   52330 => x"ffffff",
   52331 => x"ffffff",
   52332 => x"ffffff",
   52333 => x"ffffff",
   52334 => x"ffffff",
   52335 => x"ffffff",
   52336 => x"ffffff",
   52337 => x"ffffff",
   52338 => x"ffffff",
   52339 => x"ffffff",
   52340 => x"ffffff",
   52341 => x"ffffff",
   52342 => x"ffffff",
   52343 => x"ffffff",
   52344 => x"ffffff",
   52345 => x"ffffff",
   52346 => x"ffffff",
   52347 => x"ffffff",
   52348 => x"ffffff",
   52349 => x"ffffff",
   52350 => x"ffffff",
   52351 => x"ffffff",
   52352 => x"ffffff",
   52353 => x"ffffff",
   52354 => x"ffffff",
   52355 => x"ffffff",
   52356 => x"ffffff",
   52357 => x"ffffff",
   52358 => x"ffffff",
   52359 => x"ffffff",
   52360 => x"ffffff",
   52361 => x"ffffff",
   52362 => x"ffffff",
   52363 => x"ffffff",
   52364 => x"ffffff",
   52365 => x"ffffff",
   52366 => x"ffffff",
   52367 => x"ffffff",
   52368 => x"ffffff",
   52369 => x"ffffff",
   52370 => x"ffffff",
   52371 => x"ffffff",
   52372 => x"ffffff",
   52373 => x"ffffff",
   52374 => x"ffffff",
   52375 => x"ffffff",
   52376 => x"ffffff",
   52377 => x"ffffff",
   52378 => x"ffffff",
   52379 => x"ffffff",
   52380 => x"ffffff",
   52381 => x"ffffff",
   52382 => x"ffffff",
   52383 => x"ffffff",
   52384 => x"ffffff",
   52385 => x"ffffff",
   52386 => x"ffffff",
   52387 => x"ffffff",
   52388 => x"ffffff",
   52389 => x"fffa95",
   52390 => x"abffff",
   52391 => x"ffffff",
   52392 => x"ffffff",
   52393 => x"ffffff",
   52394 => x"ffffff",
   52395 => x"ffffff",
   52396 => x"ffffff",
   52397 => x"ffffff",
   52398 => x"ffffff",
   52399 => x"ffffff",
   52400 => x"ffffff",
   52401 => x"fffac3",
   52402 => x"0c30c3",
   52403 => x"0c30c3",
   52404 => x"0c30c3",
   52405 => x"0c30c3",
   52406 => x"0c30c3",
   52407 => x"0c30c3",
   52408 => x"0c30c3",
   52409 => x"0c30c3",
   52410 => x"0c30c3",
   52411 => x"0c30c3",
   52412 => x"0c30c3",
   52413 => x"082082",
   52414 => x"082082",
   52415 => x"082082",
   52416 => x"082082",
   52417 => x"082082",
   52418 => x"082082",
   52419 => x"082082",
   52420 => x"082082",
   52421 => x"082082",
   52422 => x"082082",
   52423 => x"082082",
   52424 => x"082082",
   52425 => x"082082",
   52426 => x"082082",
   52427 => x"082082",
   52428 => x"082082",
   52429 => x"082082",
   52430 => x"082082",
   52431 => x"082082",
   52432 => x"082082",
   52433 => x"082082",
   52434 => x"082082",
   52435 => x"082041",
   52436 => x"041041",
   52437 => x"041041",
   52438 => x"041041",
   52439 => x"041041",
   52440 => x"041041",
   52441 => x"041041",
   52442 => x"041041",
   52443 => x"041041",
   52444 => x"041041",
   52445 => x"041041",
   52446 => x"041041",
   52447 => x"041041",
   52448 => x"041041",
   52449 => x"041041",
   52450 => x"041041",
   52451 => x"041041",
   52452 => x"041041",
   52453 => x"041041",
   52454 => x"041041",
   52455 => x"041041",
   52456 => x"041041",
   52457 => x"041041",
   52458 => x"041000",
   52459 => x"000000",
   52460 => x"000000",
   52461 => x"000000",
   52462 => x"000000",
   52463 => x"000000",
   52464 => x"000000",
   52465 => x"000000",
   52466 => x"000000",
   52467 => x"000000",
   52468 => x"000000",
   52469 => x"00057f",
   52470 => x"ffffff",
   52471 => x"ffffff",
   52472 => x"ffffff",
   52473 => x"ffffd5",
   52474 => x"00002a",
   52475 => x"ffffff",
   52476 => x"ffffff",
   52477 => x"ffffd5",
   52478 => x"000015",
   52479 => x"ffffff",
   52480 => x"ffffff",
   52481 => x"ffffff",
   52482 => x"ffffff",
   52483 => x"ffffff",
   52484 => x"ffffff",
   52485 => x"ffffff",
   52486 => x"ffffff",
   52487 => x"ffffff",
   52488 => x"ffffff",
   52489 => x"ffffff",
   52490 => x"ffffff",
   52491 => x"ffffff",
   52492 => x"ffffff",
   52493 => x"ffffff",
   52494 => x"ffffff",
   52495 => x"ffffff",
   52496 => x"ffffff",
   52497 => x"ffffff",
   52498 => x"ffffff",
   52499 => x"ffffff",
   52500 => x"ffffff",
   52501 => x"ffffff",
   52502 => x"ffffff",
   52503 => x"ffffff",
   52504 => x"ffffff",
   52505 => x"ffffff",
   52506 => x"ffffff",
   52507 => x"ffffff",
   52508 => x"ffffff",
   52509 => x"ffffff",
   52510 => x"ffffff",
   52511 => x"ffffff",
   52512 => x"ffffff",
   52513 => x"ffffff",
   52514 => x"ffffff",
   52515 => x"ffffff",
   52516 => x"ffffff",
   52517 => x"ffffff",
   52518 => x"ffffff",
   52519 => x"ffffff",
   52520 => x"ffffff",
   52521 => x"ffffff",
   52522 => x"ffffff",
   52523 => x"ffffff",
   52524 => x"ffffff",
   52525 => x"ffffff",
   52526 => x"ffffff",
   52527 => x"ffffff",
   52528 => x"ffffff",
   52529 => x"ffffff",
   52530 => x"ffffff",
   52531 => x"ffffff",
   52532 => x"ffffff",
   52533 => x"ffffff",
   52534 => x"ffffff",
   52535 => x"ffffff",
   52536 => x"ffffff",
   52537 => x"ffffff",
   52538 => x"ffffff",
   52539 => x"ffffff",
   52540 => x"ffffff",
   52541 => x"ffffff",
   52542 => x"ffffff",
   52543 => x"ffffff",
   52544 => x"ffffff",
   52545 => x"ffffff",
   52546 => x"ffffff",
   52547 => x"ffffff",
   52548 => x"ffffff",
   52549 => x"fffa95",
   52550 => x"abffff",
   52551 => x"ffffff",
   52552 => x"ffffff",
   52553 => x"ffffff",
   52554 => x"ffffff",
   52555 => x"ffffff",
   52556 => x"ffffff",
   52557 => x"ffffff",
   52558 => x"ffffff",
   52559 => x"ffffff",
   52560 => x"ffffff",
   52561 => x"fffac3",
   52562 => x"0c30c3",
   52563 => x"0c30c3",
   52564 => x"0c30c3",
   52565 => x"0c30c3",
   52566 => x"0c30c3",
   52567 => x"0c30c3",
   52568 => x"0c30c3",
   52569 => x"0c30c3",
   52570 => x"0c30c3",
   52571 => x"0c30c3",
   52572 => x"0c30c3",
   52573 => x"082082",
   52574 => x"082082",
   52575 => x"082082",
   52576 => x"082082",
   52577 => x"082082",
   52578 => x"082082",
   52579 => x"082082",
   52580 => x"082082",
   52581 => x"082082",
   52582 => x"082082",
   52583 => x"082082",
   52584 => x"082082",
   52585 => x"082082",
   52586 => x"082082",
   52587 => x"082082",
   52588 => x"082082",
   52589 => x"082082",
   52590 => x"082082",
   52591 => x"082082",
   52592 => x"082082",
   52593 => x"082082",
   52594 => x"082082",
   52595 => x"082041",
   52596 => x"041041",
   52597 => x"041041",
   52598 => x"041041",
   52599 => x"041041",
   52600 => x"041041",
   52601 => x"041041",
   52602 => x"041041",
   52603 => x"041041",
   52604 => x"041041",
   52605 => x"041041",
   52606 => x"041041",
   52607 => x"041041",
   52608 => x"041041",
   52609 => x"041041",
   52610 => x"041041",
   52611 => x"041041",
   52612 => x"041041",
   52613 => x"041041",
   52614 => x"041041",
   52615 => x"041041",
   52616 => x"041041",
   52617 => x"041041",
   52618 => x"041000",
   52619 => x"000000",
   52620 => x"000000",
   52621 => x"000000",
   52622 => x"000000",
   52623 => x"000000",
   52624 => x"000000",
   52625 => x"000000",
   52626 => x"000000",
   52627 => x"000000",
   52628 => x"000000",
   52629 => x"00057f",
   52630 => x"ffffff",
   52631 => x"ffffff",
   52632 => x"ffffff",
   52633 => x"ffffd5",
   52634 => x"00002a",
   52635 => x"ffffff",
   52636 => x"ffffff",
   52637 => x"ffffd5",
   52638 => x"000015",
   52639 => x"ffffff",
   52640 => x"ffffff",
   52641 => x"ffffff",
   52642 => x"ffffff",
   52643 => x"ffffff",
   52644 => x"ffffff",
   52645 => x"ffffff",
   52646 => x"ffffff",
   52647 => x"ffffff",
   52648 => x"ffffff",
   52649 => x"ffffff",
   52650 => x"ffffff",
   52651 => x"ffffff",
   52652 => x"ffffff",
   52653 => x"ffffff",
   52654 => x"ffffff",
   52655 => x"ffffff",
   52656 => x"ffffff",
   52657 => x"ffffff",
   52658 => x"ffffff",
   52659 => x"ffffff",
   52660 => x"ffffff",
   52661 => x"ffffff",
   52662 => x"ffffff",
   52663 => x"ffffff",
   52664 => x"ffffff",
   52665 => x"ffffff",
   52666 => x"ffffff",
   52667 => x"ffffff",
   52668 => x"ffffff",
   52669 => x"ffffff",
   52670 => x"ffffff",
   52671 => x"ffffff",
   52672 => x"ffffff",
   52673 => x"ffffff",
   52674 => x"ffffff",
   52675 => x"ffffff",
   52676 => x"ffffff",
   52677 => x"ffffff",
   52678 => x"ffffff",
   52679 => x"ffffff",
   52680 => x"ffffff",
   52681 => x"ffffff",
   52682 => x"ffffff",
   52683 => x"ffffff",
   52684 => x"ffffff",
   52685 => x"ffffff",
   52686 => x"ffffff",
   52687 => x"ffffff",
   52688 => x"ffffff",
   52689 => x"ffffff",
   52690 => x"ffffff",
   52691 => x"ffffff",
   52692 => x"ffffff",
   52693 => x"ffffff",
   52694 => x"ffffff",
   52695 => x"ffffff",
   52696 => x"ffffff",
   52697 => x"ffffff",
   52698 => x"ffffff",
   52699 => x"ffffff",
   52700 => x"ffffff",
   52701 => x"ffffff",
   52702 => x"ffffff",
   52703 => x"ffffff",
   52704 => x"ffffff",
   52705 => x"ffffff",
   52706 => x"ffffff",
   52707 => x"ffffff",
   52708 => x"ffffff",
   52709 => x"fffa95",
   52710 => x"abffff",
   52711 => x"ffffff",
   52712 => x"ffffff",
   52713 => x"ffffff",
   52714 => x"ffffff",
   52715 => x"ffffff",
   52716 => x"ffffff",
   52717 => x"ffffff",
   52718 => x"ffffff",
   52719 => x"ffffff",
   52720 => x"ffffff",
   52721 => x"fffac3",
   52722 => x"0c30c3",
   52723 => x"0c30c3",
   52724 => x"0c30c3",
   52725 => x"0c30c3",
   52726 => x"0c30c3",
   52727 => x"0c30c3",
   52728 => x"0c30c3",
   52729 => x"0c30c3",
   52730 => x"0c30c3",
   52731 => x"0c30c3",
   52732 => x"0c30c3",
   52733 => x"082082",
   52734 => x"082082",
   52735 => x"082082",
   52736 => x"082082",
   52737 => x"082082",
   52738 => x"082082",
   52739 => x"082082",
   52740 => x"082082",
   52741 => x"082082",
   52742 => x"082082",
   52743 => x"082082",
   52744 => x"082082",
   52745 => x"082082",
   52746 => x"082082",
   52747 => x"082082",
   52748 => x"082082",
   52749 => x"082082",
   52750 => x"082082",
   52751 => x"082082",
   52752 => x"082082",
   52753 => x"082082",
   52754 => x"082082",
   52755 => x"082041",
   52756 => x"041041",
   52757 => x"041041",
   52758 => x"041041",
   52759 => x"041041",
   52760 => x"041041",
   52761 => x"041041",
   52762 => x"041041",
   52763 => x"041041",
   52764 => x"041041",
   52765 => x"041041",
   52766 => x"041041",
   52767 => x"041041",
   52768 => x"041041",
   52769 => x"041041",
   52770 => x"041041",
   52771 => x"041041",
   52772 => x"041041",
   52773 => x"041041",
   52774 => x"041041",
   52775 => x"041041",
   52776 => x"041041",
   52777 => x"041041",
   52778 => x"041000",
   52779 => x"000000",
   52780 => x"000000",
   52781 => x"000000",
   52782 => x"000000",
   52783 => x"000000",
   52784 => x"000000",
   52785 => x"000000",
   52786 => x"000000",
   52787 => x"000000",
   52788 => x"000000",
   52789 => x"00057f",
   52790 => x"ffffff",
   52791 => x"ffffff",
   52792 => x"ffffff",
   52793 => x"ffffd5",
   52794 => x"00002a",
   52795 => x"ffffff",
   52796 => x"ffffff",
   52797 => x"ffffd5",
   52798 => x"00002a",
   52799 => x"ffffff",
   52800 => x"ffffff",
   52801 => x"ffffff",
   52802 => x"ffffff",
   52803 => x"ffffff",
   52804 => x"ffffff",
   52805 => x"ffffff",
   52806 => x"ffffff",
   52807 => x"ffffff",
   52808 => x"ffffff",
   52809 => x"ffffff",
   52810 => x"ffffff",
   52811 => x"ffffff",
   52812 => x"ffffff",
   52813 => x"ffffff",
   52814 => x"ffffff",
   52815 => x"ffffff",
   52816 => x"ffffff",
   52817 => x"ffffff",
   52818 => x"ffffff",
   52819 => x"ffffff",
   52820 => x"ffffff",
   52821 => x"ffffff",
   52822 => x"ffffff",
   52823 => x"ffffff",
   52824 => x"ffffff",
   52825 => x"ffffff",
   52826 => x"ffffff",
   52827 => x"ffffff",
   52828 => x"ffffff",
   52829 => x"ffffff",
   52830 => x"ffffff",
   52831 => x"ffffff",
   52832 => x"ffffff",
   52833 => x"ffffff",
   52834 => x"ffffff",
   52835 => x"ffffff",
   52836 => x"ffffff",
   52837 => x"ffffff",
   52838 => x"ffffff",
   52839 => x"ffffff",
   52840 => x"ffffff",
   52841 => x"ffffff",
   52842 => x"ffffff",
   52843 => x"ffffff",
   52844 => x"ffffff",
   52845 => x"ffffff",
   52846 => x"ffffff",
   52847 => x"ffffff",
   52848 => x"ffffff",
   52849 => x"ffffff",
   52850 => x"ffffff",
   52851 => x"ffffff",
   52852 => x"ffffff",
   52853 => x"ffffff",
   52854 => x"ffffff",
   52855 => x"ffffff",
   52856 => x"ffffff",
   52857 => x"ffffff",
   52858 => x"ffffff",
   52859 => x"ffffff",
   52860 => x"ffffff",
   52861 => x"ffffff",
   52862 => x"ffffff",
   52863 => x"ffffff",
   52864 => x"ffffff",
   52865 => x"ffffff",
   52866 => x"ffffff",
   52867 => x"ffffff",
   52868 => x"ffffff",
   52869 => x"fffa95",
   52870 => x"abffff",
   52871 => x"ffffff",
   52872 => x"ffffff",
   52873 => x"ffffff",
   52874 => x"ffffff",
   52875 => x"ffffff",
   52876 => x"ffffff",
   52877 => x"ffffff",
   52878 => x"ffffff",
   52879 => x"ffffff",
   52880 => x"ffffff",
   52881 => x"fffac3",
   52882 => x"0c30c3",
   52883 => x"0c30c3",
   52884 => x"0c30c3",
   52885 => x"0c30c3",
   52886 => x"0c30c3",
   52887 => x"0c30c3",
   52888 => x"0c30c3",
   52889 => x"0c30c3",
   52890 => x"0c30c3",
   52891 => x"0c30c3",
   52892 => x"0c30c3",
   52893 => x"082082",
   52894 => x"082082",
   52895 => x"082082",
   52896 => x"082082",
   52897 => x"082082",
   52898 => x"082082",
   52899 => x"082082",
   52900 => x"082082",
   52901 => x"082082",
   52902 => x"082082",
   52903 => x"082082",
   52904 => x"082082",
   52905 => x"082082",
   52906 => x"082082",
   52907 => x"082082",
   52908 => x"082082",
   52909 => x"082082",
   52910 => x"082082",
   52911 => x"082082",
   52912 => x"082082",
   52913 => x"082082",
   52914 => x"082082",
   52915 => x"082041",
   52916 => x"041041",
   52917 => x"041041",
   52918 => x"041041",
   52919 => x"041041",
   52920 => x"041041",
   52921 => x"041041",
   52922 => x"041041",
   52923 => x"041041",
   52924 => x"041041",
   52925 => x"041041",
   52926 => x"041041",
   52927 => x"041041",
   52928 => x"041041",
   52929 => x"041041",
   52930 => x"041041",
   52931 => x"041041",
   52932 => x"041041",
   52933 => x"041041",
   52934 => x"041041",
   52935 => x"041041",
   52936 => x"041041",
   52937 => x"041041",
   52938 => x"041000",
   52939 => x"000000",
   52940 => x"000000",
   52941 => x"000000",
   52942 => x"000000",
   52943 => x"000000",
   52944 => x"000000",
   52945 => x"000000",
   52946 => x"000000",
   52947 => x"000000",
   52948 => x"000000",
   52949 => x"00057f",
   52950 => x"ffffff",
   52951 => x"ffffff",
   52952 => x"ffffff",
   52953 => x"ffffd5",
   52954 => x"00002a",
   52955 => x"ffffff",
   52956 => x"ffffff",
   52957 => x"fffa95",
   52958 => x"00002a",
   52959 => x"ffffff",
   52960 => x"ffffff",
   52961 => x"ffffff",
   52962 => x"ffffff",
   52963 => x"ffffff",
   52964 => x"ffffff",
   52965 => x"ffffff",
   52966 => x"ffffff",
   52967 => x"ffffff",
   52968 => x"ffffff",
   52969 => x"ffffff",
   52970 => x"ffffff",
   52971 => x"ffffff",
   52972 => x"ffffff",
   52973 => x"ffffff",
   52974 => x"ffffff",
   52975 => x"ffffff",
   52976 => x"ffffff",
   52977 => x"ffffff",
   52978 => x"ffffff",
   52979 => x"ffffff",
   52980 => x"ffffff",
   52981 => x"ffffff",
   52982 => x"ffffff",
   52983 => x"ffffff",
   52984 => x"ffffff",
   52985 => x"ffffff",
   52986 => x"ffffff",
   52987 => x"ffffff",
   52988 => x"ffffff",
   52989 => x"ffffff",
   52990 => x"ffffff",
   52991 => x"ffffff",
   52992 => x"ffffff",
   52993 => x"ffffff",
   52994 => x"ffffff",
   52995 => x"ffffff",
   52996 => x"ffffff",
   52997 => x"ffffff",
   52998 => x"ffffff",
   52999 => x"ffffff",
   53000 => x"ffffff",
   53001 => x"ffffff",
   53002 => x"ffffff",
   53003 => x"ffffff",
   53004 => x"ffffff",
   53005 => x"ffffff",
   53006 => x"ffffff",
   53007 => x"ffffff",
   53008 => x"ffffff",
   53009 => x"ffffff",
   53010 => x"ffffff",
   53011 => x"ffffff",
   53012 => x"ffffff",
   53013 => x"ffffff",
   53014 => x"ffffff",
   53015 => x"ffffff",
   53016 => x"ffffff",
   53017 => x"ffffff",
   53018 => x"ffffff",
   53019 => x"ffffff",
   53020 => x"ffffff",
   53021 => x"ffffff",
   53022 => x"ffffff",
   53023 => x"ffffff",
   53024 => x"ffffff",
   53025 => x"ffffff",
   53026 => x"ffffff",
   53027 => x"ffffff",
   53028 => x"ffffff",
   53029 => x"fffa95",
   53030 => x"abffff",
   53031 => x"ffffff",
   53032 => x"ffffff",
   53033 => x"ffffff",
   53034 => x"ffffff",
   53035 => x"ffffff",
   53036 => x"ffffff",
   53037 => x"ffffff",
   53038 => x"ffffff",
   53039 => x"ffffff",
   53040 => x"ffffff",
   53041 => x"fffac3",
   53042 => x"0c30c3",
   53043 => x"0c30c3",
   53044 => x"0c30c3",
   53045 => x"0c30c3",
   53046 => x"0c30c3",
   53047 => x"0c30c3",
   53048 => x"0c30c3",
   53049 => x"0c30c3",
   53050 => x"0c30c3",
   53051 => x"0c30c3",
   53052 => x"0c30c3",
   53053 => x"082082",
   53054 => x"082082",
   53055 => x"082082",
   53056 => x"082082",
   53057 => x"082082",
   53058 => x"082082",
   53059 => x"082082",
   53060 => x"082082",
   53061 => x"082082",
   53062 => x"082082",
   53063 => x"082082",
   53064 => x"082082",
   53065 => x"082082",
   53066 => x"082082",
   53067 => x"082082",
   53068 => x"082082",
   53069 => x"082082",
   53070 => x"082082",
   53071 => x"082082",
   53072 => x"082082",
   53073 => x"082082",
   53074 => x"082082",
   53075 => x"082041",
   53076 => x"041041",
   53077 => x"041041",
   53078 => x"041041",
   53079 => x"041041",
   53080 => x"041041",
   53081 => x"041041",
   53082 => x"041041",
   53083 => x"041041",
   53084 => x"041041",
   53085 => x"041041",
   53086 => x"041041",
   53087 => x"041041",
   53088 => x"041041",
   53089 => x"041041",
   53090 => x"041041",
   53091 => x"041041",
   53092 => x"041041",
   53093 => x"041041",
   53094 => x"041041",
   53095 => x"041041",
   53096 => x"041041",
   53097 => x"041041",
   53098 => x"041000",
   53099 => x"000000",
   53100 => x"000000",
   53101 => x"000000",
   53102 => x"000000",
   53103 => x"000000",
   53104 => x"000000",
   53105 => x"000000",
   53106 => x"000000",
   53107 => x"000000",
   53108 => x"000000",
   53109 => x"00057f",
   53110 => x"ffffff",
   53111 => x"ffffff",
   53112 => x"ffffff",
   53113 => x"ffffd5",
   53114 => x"00002a",
   53115 => x"ffffff",
   53116 => x"ffffff",
   53117 => x"fff540",
   53118 => x"00057f",
   53119 => x"ffffff",
   53120 => x"ffffff",
   53121 => x"ffffff",
   53122 => x"ffffff",
   53123 => x"ffffff",
   53124 => x"ffffff",
   53125 => x"ffffff",
   53126 => x"ffffff",
   53127 => x"ffffff",
   53128 => x"ffffff",
   53129 => x"ffffff",
   53130 => x"ffffff",
   53131 => x"ffffff",
   53132 => x"ffffff",
   53133 => x"ffffff",
   53134 => x"ffffff",
   53135 => x"ffffff",
   53136 => x"ffffff",
   53137 => x"ffffff",
   53138 => x"ffffff",
   53139 => x"ffffff",
   53140 => x"ffffff",
   53141 => x"ffffff",
   53142 => x"ffffff",
   53143 => x"ffffff",
   53144 => x"ffffff",
   53145 => x"ffffff",
   53146 => x"ffffff",
   53147 => x"ffffff",
   53148 => x"ffffff",
   53149 => x"ffffff",
   53150 => x"ffffff",
   53151 => x"ffffff",
   53152 => x"ffffff",
   53153 => x"ffffff",
   53154 => x"ffffff",
   53155 => x"ffffff",
   53156 => x"ffffff",
   53157 => x"ffffff",
   53158 => x"ffffff",
   53159 => x"ffffff",
   53160 => x"ffffff",
   53161 => x"ffffff",
   53162 => x"ffffff",
   53163 => x"ffffff",
   53164 => x"ffffff",
   53165 => x"ffffff",
   53166 => x"ffffff",
   53167 => x"ffffff",
   53168 => x"ffffff",
   53169 => x"ffffff",
   53170 => x"ffffff",
   53171 => x"ffffff",
   53172 => x"ffffff",
   53173 => x"ffffff",
   53174 => x"ffffff",
   53175 => x"ffffff",
   53176 => x"ffffff",
   53177 => x"ffffff",
   53178 => x"ffffff",
   53179 => x"ffffff",
   53180 => x"ffffff",
   53181 => x"ffffff",
   53182 => x"ffffff",
   53183 => x"ffffff",
   53184 => x"ffffff",
   53185 => x"ffffff",
   53186 => x"ffffff",
   53187 => x"ffffff",
   53188 => x"ffffff",
   53189 => x"fffa95",
   53190 => x"abffff",
   53191 => x"ffffff",
   53192 => x"ffffff",
   53193 => x"ffffff",
   53194 => x"ffffff",
   53195 => x"ffffff",
   53196 => x"ffffff",
   53197 => x"ffffff",
   53198 => x"ffffff",
   53199 => x"ffffff",
   53200 => x"ffffff",
   53201 => x"fffac3",
   53202 => x"0c30c3",
   53203 => x"0c30c3",
   53204 => x"0c30c3",
   53205 => x"0c30c3",
   53206 => x"0c30c3",
   53207 => x"0c30c3",
   53208 => x"0c30c3",
   53209 => x"0c30c3",
   53210 => x"0c30c3",
   53211 => x"0c30c3",
   53212 => x"0c30c3",
   53213 => x"082082",
   53214 => x"082082",
   53215 => x"082082",
   53216 => x"082082",
   53217 => x"082082",
   53218 => x"082082",
   53219 => x"082082",
   53220 => x"082082",
   53221 => x"082082",
   53222 => x"082082",
   53223 => x"082082",
   53224 => x"082082",
   53225 => x"082082",
   53226 => x"082082",
   53227 => x"082082",
   53228 => x"082082",
   53229 => x"082082",
   53230 => x"082082",
   53231 => x"082082",
   53232 => x"082082",
   53233 => x"082082",
   53234 => x"082082",
   53235 => x"082041",
   53236 => x"041041",
   53237 => x"041041",
   53238 => x"041041",
   53239 => x"041041",
   53240 => x"041041",
   53241 => x"041041",
   53242 => x"041041",
   53243 => x"041041",
   53244 => x"041041",
   53245 => x"041041",
   53246 => x"041041",
   53247 => x"041041",
   53248 => x"041041",
   53249 => x"041041",
   53250 => x"041041",
   53251 => x"041041",
   53252 => x"041041",
   53253 => x"041041",
   53254 => x"041041",
   53255 => x"041041",
   53256 => x"041041",
   53257 => x"041041",
   53258 => x"041000",
   53259 => x"000000",
   53260 => x"000000",
   53261 => x"000000",
   53262 => x"000000",
   53263 => x"000000",
   53264 => x"000000",
   53265 => x"000000",
   53266 => x"000000",
   53267 => x"000000",
   53268 => x"000000",
   53269 => x"00057f",
   53270 => x"ffffff",
   53271 => x"ffffff",
   53272 => x"ffffff",
   53273 => x"ffffd5",
   53274 => x"00002a",
   53275 => x"ffffff",
   53276 => x"ffffea",
   53277 => x"a95000",
   53278 => x"000abf",
   53279 => x"ffffff",
   53280 => x"ffffff",
   53281 => x"ffffff",
   53282 => x"ffffff",
   53283 => x"ffffff",
   53284 => x"ffffff",
   53285 => x"ffffff",
   53286 => x"ffffff",
   53287 => x"ffffff",
   53288 => x"ffffff",
   53289 => x"ffffff",
   53290 => x"ffffff",
   53291 => x"ffffff",
   53292 => x"ffffff",
   53293 => x"ffffff",
   53294 => x"ffffff",
   53295 => x"ffffff",
   53296 => x"ffffff",
   53297 => x"ffffff",
   53298 => x"ffffff",
   53299 => x"ffffff",
   53300 => x"ffffff",
   53301 => x"ffffff",
   53302 => x"ffffff",
   53303 => x"ffffff",
   53304 => x"ffffff",
   53305 => x"ffffff",
   53306 => x"ffffff",
   53307 => x"ffffff",
   53308 => x"ffffff",
   53309 => x"ffffff",
   53310 => x"ffffff",
   53311 => x"ffffff",
   53312 => x"ffffff",
   53313 => x"ffffff",
   53314 => x"ffffff",
   53315 => x"ffffff",
   53316 => x"ffffff",
   53317 => x"ffffff",
   53318 => x"ffffff",
   53319 => x"ffffff",
   53320 => x"ffffff",
   53321 => x"ffffff",
   53322 => x"ffffff",
   53323 => x"ffffff",
   53324 => x"ffffff",
   53325 => x"ffffff",
   53326 => x"ffffff",
   53327 => x"ffffff",
   53328 => x"ffffff",
   53329 => x"ffffff",
   53330 => x"ffffff",
   53331 => x"ffffff",
   53332 => x"ffffff",
   53333 => x"ffffff",
   53334 => x"ffffff",
   53335 => x"ffffff",
   53336 => x"ffffff",
   53337 => x"ffffff",
   53338 => x"ffffff",
   53339 => x"ffffff",
   53340 => x"ffffff",
   53341 => x"ffffff",
   53342 => x"ffffff",
   53343 => x"ffffff",
   53344 => x"ffffff",
   53345 => x"ffffff",
   53346 => x"ffffff",
   53347 => x"ffffff",
   53348 => x"ffffff",
   53349 => x"fffa95",
   53350 => x"abffff",
   53351 => x"ffffff",
   53352 => x"ffffff",
   53353 => x"ffffff",
   53354 => x"ffffff",
   53355 => x"ffffff",
   53356 => x"ffffff",
   53357 => x"ffffff",
   53358 => x"ffffff",
   53359 => x"ffffff",
   53360 => x"ffffff",
   53361 => x"fffac3",
   53362 => x"0c30c3",
   53363 => x"0c30c3",
   53364 => x"0c30c3",
   53365 => x"0c30c3",
   53366 => x"0c30c3",
   53367 => x"0c30c3",
   53368 => x"0c30c3",
   53369 => x"0c30c3",
   53370 => x"0c30c3",
   53371 => x"0c30c3",
   53372 => x"0c30c3",
   53373 => x"082082",
   53374 => x"082082",
   53375 => x"082082",
   53376 => x"082082",
   53377 => x"082082",
   53378 => x"082082",
   53379 => x"082082",
   53380 => x"082082",
   53381 => x"082082",
   53382 => x"082082",
   53383 => x"082082",
   53384 => x"082082",
   53385 => x"082082",
   53386 => x"082082",
   53387 => x"082082",
   53388 => x"082082",
   53389 => x"082082",
   53390 => x"082082",
   53391 => x"082082",
   53392 => x"082082",
   53393 => x"082082",
   53394 => x"082082",
   53395 => x"082041",
   53396 => x"041041",
   53397 => x"041041",
   53398 => x"041041",
   53399 => x"041041",
   53400 => x"041041",
   53401 => x"041041",
   53402 => x"041041",
   53403 => x"041041",
   53404 => x"041041",
   53405 => x"041041",
   53406 => x"041041",
   53407 => x"041041",
   53408 => x"041041",
   53409 => x"041041",
   53410 => x"041041",
   53411 => x"041041",
   53412 => x"041041",
   53413 => x"041041",
   53414 => x"041041",
   53415 => x"041041",
   53416 => x"041041",
   53417 => x"041041",
   53418 => x"041000",
   53419 => x"000000",
   53420 => x"000000",
   53421 => x"000000",
   53422 => x"000000",
   53423 => x"000000",
   53424 => x"000000",
   53425 => x"000000",
   53426 => x"000000",
   53427 => x"000000",
   53428 => x"000000",
   53429 => x"00057f",
   53430 => x"ffffff",
   53431 => x"ffffff",
   53432 => x"ffffff",
   53433 => x"ffffd5",
   53434 => x"000015",
   53435 => x"555555",
   53436 => x"555555",
   53437 => x"000000",
   53438 => x"56afff",
   53439 => x"ffffff",
   53440 => x"ffffff",
   53441 => x"ffffff",
   53442 => x"ffffff",
   53443 => x"ffffff",
   53444 => x"ffffff",
   53445 => x"ffffff",
   53446 => x"ffffff",
   53447 => x"ffffff",
   53448 => x"ffffff",
   53449 => x"ffffff",
   53450 => x"ffffff",
   53451 => x"ffffff",
   53452 => x"ffffff",
   53453 => x"ffffff",
   53454 => x"ffffff",
   53455 => x"ffffff",
   53456 => x"ffffff",
   53457 => x"ffffff",
   53458 => x"ffffff",
   53459 => x"ffffff",
   53460 => x"ffffff",
   53461 => x"ffffff",
   53462 => x"ffffff",
   53463 => x"ffffff",
   53464 => x"ffffff",
   53465 => x"ffffff",
   53466 => x"ffffff",
   53467 => x"ffffff",
   53468 => x"ffffff",
   53469 => x"ffffff",
   53470 => x"ffffff",
   53471 => x"ffffff",
   53472 => x"ffffff",
   53473 => x"ffffff",
   53474 => x"ffffff",
   53475 => x"ffffff",
   53476 => x"ffffff",
   53477 => x"ffffff",
   53478 => x"ffffff",
   53479 => x"ffffff",
   53480 => x"ffffff",
   53481 => x"ffffff",
   53482 => x"ffffff",
   53483 => x"ffffff",
   53484 => x"ffffff",
   53485 => x"ffffff",
   53486 => x"ffffff",
   53487 => x"ffffff",
   53488 => x"ffffff",
   53489 => x"ffffff",
   53490 => x"ffffff",
   53491 => x"ffffff",
   53492 => x"ffffff",
   53493 => x"ffffff",
   53494 => x"ffffff",
   53495 => x"ffffff",
   53496 => x"ffffff",
   53497 => x"ffffff",
   53498 => x"ffffff",
   53499 => x"ffffff",
   53500 => x"ffffff",
   53501 => x"ffffff",
   53502 => x"ffffff",
   53503 => x"ffffff",
   53504 => x"ffffff",
   53505 => x"ffffff",
   53506 => x"ffffff",
   53507 => x"ffffff",
   53508 => x"ffffff",
   53509 => x"fffa95",
   53510 => x"abffff",
   53511 => x"ffffff",
   53512 => x"ffffff",
   53513 => x"ffffff",
   53514 => x"ffffff",
   53515 => x"ffffff",
   53516 => x"ffffff",
   53517 => x"ffffff",
   53518 => x"ffffff",
   53519 => x"ffffff",
   53520 => x"ffffff",
   53521 => x"fffac3",
   53522 => x"0c30c3",
   53523 => x"0c30c3",
   53524 => x"0c30c3",
   53525 => x"0c30c3",
   53526 => x"0c30c3",
   53527 => x"0c30c3",
   53528 => x"0c30c3",
   53529 => x"0c30c3",
   53530 => x"0c30c3",
   53531 => x"0c30c3",
   53532 => x"0c30c3",
   53533 => x"082082",
   53534 => x"082082",
   53535 => x"082082",
   53536 => x"082082",
   53537 => x"082082",
   53538 => x"082082",
   53539 => x"082082",
   53540 => x"082082",
   53541 => x"082082",
   53542 => x"082082",
   53543 => x"082082",
   53544 => x"082082",
   53545 => x"082082",
   53546 => x"082082",
   53547 => x"082082",
   53548 => x"082082",
   53549 => x"082082",
   53550 => x"082082",
   53551 => x"082082",
   53552 => x"082082",
   53553 => x"082082",
   53554 => x"082082",
   53555 => x"082041",
   53556 => x"041041",
   53557 => x"041041",
   53558 => x"041041",
   53559 => x"041041",
   53560 => x"041041",
   53561 => x"041041",
   53562 => x"041041",
   53563 => x"041041",
   53564 => x"041041",
   53565 => x"041041",
   53566 => x"041041",
   53567 => x"041041",
   53568 => x"041041",
   53569 => x"041041",
   53570 => x"041041",
   53571 => x"041041",
   53572 => x"041041",
   53573 => x"041041",
   53574 => x"041041",
   53575 => x"041041",
   53576 => x"041041",
   53577 => x"041041",
   53578 => x"041000",
   53579 => x"000000",
   53580 => x"000000",
   53581 => x"000000",
   53582 => x"000000",
   53583 => x"000000",
   53584 => x"000000",
   53585 => x"000000",
   53586 => x"000000",
   53587 => x"000000",
   53588 => x"000000",
   53589 => x"00057f",
   53590 => x"ffffff",
   53591 => x"ffffff",
   53592 => x"ffffff",
   53593 => x"ffffd5",
   53594 => x"000000",
   53595 => x"000000",
   53596 => x"000000",
   53597 => x"000015",
   53598 => x"abffff",
   53599 => x"ffffff",
   53600 => x"ffffff",
   53601 => x"ffffff",
   53602 => x"ffffff",
   53603 => x"ffffff",
   53604 => x"ffffff",
   53605 => x"ffffff",
   53606 => x"ffffff",
   53607 => x"ffffff",
   53608 => x"ffffff",
   53609 => x"ffffff",
   53610 => x"ffffff",
   53611 => x"ffffff",
   53612 => x"ffffff",
   53613 => x"ffffff",
   53614 => x"ffffff",
   53615 => x"ffffff",
   53616 => x"ffffff",
   53617 => x"ffffff",
   53618 => x"ffffff",
   53619 => x"ffffff",
   53620 => x"ffffff",
   53621 => x"ffffff",
   53622 => x"ffffff",
   53623 => x"ffffff",
   53624 => x"ffffff",
   53625 => x"ffffff",
   53626 => x"ffffff",
   53627 => x"ffffff",
   53628 => x"ffffff",
   53629 => x"ffffff",
   53630 => x"ffffff",
   53631 => x"ffffff",
   53632 => x"ffffff",
   53633 => x"ffffff",
   53634 => x"ffffff",
   53635 => x"ffffff",
   53636 => x"ffffff",
   53637 => x"ffffff",
   53638 => x"ffffff",
   53639 => x"ffffff",
   53640 => x"ffffff",
   53641 => x"ffffff",
   53642 => x"ffffff",
   53643 => x"ffffff",
   53644 => x"ffffff",
   53645 => x"ffffff",
   53646 => x"ffffff",
   53647 => x"ffffff",
   53648 => x"ffffff",
   53649 => x"ffffff",
   53650 => x"ffffff",
   53651 => x"ffffff",
   53652 => x"ffffff",
   53653 => x"ffffff",
   53654 => x"ffffff",
   53655 => x"ffffff",
   53656 => x"ffffff",
   53657 => x"ffffff",
   53658 => x"ffffff",
   53659 => x"ffffff",
   53660 => x"ffffff",
   53661 => x"ffffff",
   53662 => x"ffffff",
   53663 => x"ffffff",
   53664 => x"ffffff",
   53665 => x"ffffff",
   53666 => x"ffffff",
   53667 => x"ffffff",
   53668 => x"ffffff",
   53669 => x"fffa95",
   53670 => x"abffff",
   53671 => x"ffffff",
   53672 => x"ffffff",
   53673 => x"ffffff",
   53674 => x"ffffff",
   53675 => x"ffffff",
   53676 => x"ffffff",
   53677 => x"ffffff",
   53678 => x"ffffff",
   53679 => x"ffffff",
   53680 => x"ffffff",
   53681 => x"fffac3",
   53682 => x"0c30c3",
   53683 => x"0c30c3",
   53684 => x"0c30c3",
   53685 => x"0c30c3",
   53686 => x"0c30c3",
   53687 => x"0c30c3",
   53688 => x"0c30c3",
   53689 => x"0c30c3",
   53690 => x"0c30c3",
   53691 => x"0c30c3",
   53692 => x"0c30c3",
   53693 => x"082082",
   53694 => x"082082",
   53695 => x"082082",
   53696 => x"082082",
   53697 => x"082082",
   53698 => x"082082",
   53699 => x"082082",
   53700 => x"082082",
   53701 => x"082082",
   53702 => x"082082",
   53703 => x"082082",
   53704 => x"082082",
   53705 => x"082082",
   53706 => x"082082",
   53707 => x"082082",
   53708 => x"082082",
   53709 => x"082082",
   53710 => x"082082",
   53711 => x"082082",
   53712 => x"082082",
   53713 => x"082082",
   53714 => x"082082",
   53715 => x"082041",
   53716 => x"041041",
   53717 => x"041041",
   53718 => x"041041",
   53719 => x"041041",
   53720 => x"041041",
   53721 => x"041041",
   53722 => x"041041",
   53723 => x"041041",
   53724 => x"041041",
   53725 => x"041041",
   53726 => x"041041",
   53727 => x"041041",
   53728 => x"041041",
   53729 => x"041041",
   53730 => x"041041",
   53731 => x"041041",
   53732 => x"041041",
   53733 => x"041041",
   53734 => x"041041",
   53735 => x"041041",
   53736 => x"041041",
   53737 => x"041041",
   53738 => x"041000",
   53739 => x"000000",
   53740 => x"000000",
   53741 => x"000000",
   53742 => x"000000",
   53743 => x"000000",
   53744 => x"000000",
   53745 => x"000000",
   53746 => x"000000",
   53747 => x"000000",
   53748 => x"000000",
   53749 => x"00057f",
   53750 => x"ffffff",
   53751 => x"ffffff",
   53752 => x"ffffff",
   53753 => x"ffffd5",
   53754 => x"000000",
   53755 => x"000000",
   53756 => x"000000",
   53757 => x"000015",
   53758 => x"abffff",
   53759 => x"ffffff",
   53760 => x"ffffff",
   53761 => x"ffffff",
   53762 => x"ffffff",
   53763 => x"ffffff",
   53764 => x"ffffff",
   53765 => x"ffffff",
   53766 => x"ffffff",
   53767 => x"ffffff",
   53768 => x"ffffff",
   53769 => x"ffffff",
   53770 => x"ffffff",
   53771 => x"ffffff",
   53772 => x"ffffff",
   53773 => x"ffffff",
   53774 => x"ffffff",
   53775 => x"ffffff",
   53776 => x"ffffff",
   53777 => x"ffffff",
   53778 => x"ffffff",
   53779 => x"ffffff",
   53780 => x"ffffff",
   53781 => x"ffffff",
   53782 => x"ffffff",
   53783 => x"ffffff",
   53784 => x"ffffff",
   53785 => x"ffffff",
   53786 => x"ffffff",
   53787 => x"ffffff",
   53788 => x"ffffff",
   53789 => x"ffffff",
   53790 => x"ffffff",
   53791 => x"ffffff",
   53792 => x"ffffff",
   53793 => x"ffffff",
   53794 => x"ffffff",
   53795 => x"ffffff",
   53796 => x"ffffff",
   53797 => x"ffffff",
   53798 => x"ffffff",
   53799 => x"ffffff",
   53800 => x"ffffff",
   53801 => x"ffffff",
   53802 => x"ffffff",
   53803 => x"ffffff",
   53804 => x"ffffff",
   53805 => x"ffffff",
   53806 => x"ffffff",
   53807 => x"ffffff",
   53808 => x"ffffff",
   53809 => x"ffffff",
   53810 => x"ffffff",
   53811 => x"ffffff",
   53812 => x"ffffff",
   53813 => x"ffffff",
   53814 => x"ffffff",
   53815 => x"ffffff",
   53816 => x"ffffff",
   53817 => x"ffffff",
   53818 => x"ffffff",
   53819 => x"ffffff",
   53820 => x"ffffff",
   53821 => x"ffffff",
   53822 => x"ffffff",
   53823 => x"ffffff",
   53824 => x"ffffff",
   53825 => x"ffffff",
   53826 => x"ffffff",
   53827 => x"ffffff",
   53828 => x"ffffff",
   53829 => x"fffa95",
   53830 => x"abffff",
   53831 => x"ffffff",
   53832 => x"ffffff",
   53833 => x"ffffff",
   53834 => x"ffffff",
   53835 => x"ffffff",
   53836 => x"ffffff",
   53837 => x"ffffff",
   53838 => x"ffffff",
   53839 => x"ffffff",
   53840 => x"ffffff",
   53841 => x"fffac3",
   53842 => x"0c30c3",
   53843 => x"0c30c3",
   53844 => x"0c30c3",
   53845 => x"0c30c3",
   53846 => x"0c30c3",
   53847 => x"0c30c3",
   53848 => x"0c30c3",
   53849 => x"0c30c3",
   53850 => x"0c30c3",
   53851 => x"0c30c3",
   53852 => x"0c30c3",
   53853 => x"082082",
   53854 => x"082082",
   53855 => x"082082",
   53856 => x"082082",
   53857 => x"082082",
   53858 => x"082082",
   53859 => x"082082",
   53860 => x"082082",
   53861 => x"082082",
   53862 => x"082082",
   53863 => x"082082",
   53864 => x"082082",
   53865 => x"082082",
   53866 => x"082082",
   53867 => x"082082",
   53868 => x"082082",
   53869 => x"082082",
   53870 => x"082082",
   53871 => x"082082",
   53872 => x"082082",
   53873 => x"082082",
   53874 => x"082082",
   53875 => x"082041",
   53876 => x"041041",
   53877 => x"041041",
   53878 => x"041041",
   53879 => x"041041",
   53880 => x"041041",
   53881 => x"041041",
   53882 => x"041041",
   53883 => x"041041",
   53884 => x"041041",
   53885 => x"041041",
   53886 => x"041041",
   53887 => x"041041",
   53888 => x"041041",
   53889 => x"041041",
   53890 => x"041041",
   53891 => x"041041",
   53892 => x"041041",
   53893 => x"041041",
   53894 => x"041041",
   53895 => x"041041",
   53896 => x"041041",
   53897 => x"041041",
   53898 => x"041000",
   53899 => x"000000",
   53900 => x"000000",
   53901 => x"000000",
   53902 => x"000000",
   53903 => x"000000",
   53904 => x"000000",
   53905 => x"000000",
   53906 => x"000000",
   53907 => x"000000",
   53908 => x"000000",
   53909 => x"00057f",
   53910 => x"ffffff",
   53911 => x"ffffff",
   53912 => x"ffffff",
   53913 => x"ffffd5",
   53914 => x"000015",
   53915 => x"555555",
   53916 => x"555555",
   53917 => x"000000",
   53918 => x"015abf",
   53919 => x"ffffff",
   53920 => x"ffffff",
   53921 => x"ffffff",
   53922 => x"ffffff",
   53923 => x"ffffff",
   53924 => x"ffffff",
   53925 => x"ffffff",
   53926 => x"ffffff",
   53927 => x"ffffff",
   53928 => x"ffffff",
   53929 => x"ffffff",
   53930 => x"ffffff",
   53931 => x"ffffff",
   53932 => x"ffffff",
   53933 => x"ffffff",
   53934 => x"ffffff",
   53935 => x"ffffff",
   53936 => x"ffffff",
   53937 => x"ffffff",
   53938 => x"ffffff",
   53939 => x"ffffff",
   53940 => x"ffffff",
   53941 => x"ffffff",
   53942 => x"ffffff",
   53943 => x"ffffff",
   53944 => x"ffffff",
   53945 => x"ffffff",
   53946 => x"ffffff",
   53947 => x"ffffff",
   53948 => x"ffffff",
   53949 => x"ffffff",
   53950 => x"ffffff",
   53951 => x"ffffff",
   53952 => x"ffffff",
   53953 => x"ffffff",
   53954 => x"ffffff",
   53955 => x"ffffff",
   53956 => x"ffffff",
   53957 => x"ffffff",
   53958 => x"ffffff",
   53959 => x"ffffff",
   53960 => x"ffffff",
   53961 => x"ffffff",
   53962 => x"ffffff",
   53963 => x"ffffff",
   53964 => x"ffffff",
   53965 => x"ffffff",
   53966 => x"ffffff",
   53967 => x"ffffff",
   53968 => x"ffffff",
   53969 => x"ffffff",
   53970 => x"ffffff",
   53971 => x"ffffff",
   53972 => x"ffffff",
   53973 => x"ffffff",
   53974 => x"ffffff",
   53975 => x"ffffff",
   53976 => x"ffffff",
   53977 => x"ffffff",
   53978 => x"ffffff",
   53979 => x"ffffff",
   53980 => x"ffffff",
   53981 => x"ffffff",
   53982 => x"ffffff",
   53983 => x"ffffff",
   53984 => x"ffffff",
   53985 => x"ffffff",
   53986 => x"ffffff",
   53987 => x"ffffff",
   53988 => x"ffffff",
   53989 => x"fffa95",
   53990 => x"abffff",
   53991 => x"ffffff",
   53992 => x"ffffff",
   53993 => x"ffffff",
   53994 => x"ffffff",
   53995 => x"ffffff",
   53996 => x"ffffff",
   53997 => x"ffffff",
   53998 => x"ffffff",
   53999 => x"ffffff",
   54000 => x"ffffff",
   54001 => x"fffac3",
   54002 => x"0c30c3",
   54003 => x"0c30c3",
   54004 => x"0c30c3",
   54005 => x"0c30c3",
   54006 => x"0c30c3",
   54007 => x"0c30c3",
   54008 => x"0c30c3",
   54009 => x"0c30c3",
   54010 => x"0c30c3",
   54011 => x"0c30c3",
   54012 => x"0c30c3",
   54013 => x"082082",
   54014 => x"082082",
   54015 => x"082082",
   54016 => x"082082",
   54017 => x"082082",
   54018 => x"082082",
   54019 => x"082082",
   54020 => x"082082",
   54021 => x"082082",
   54022 => x"082082",
   54023 => x"082082",
   54024 => x"082082",
   54025 => x"082082",
   54026 => x"082082",
   54027 => x"082082",
   54028 => x"082082",
   54029 => x"082082",
   54030 => x"082082",
   54031 => x"082082",
   54032 => x"082082",
   54033 => x"082082",
   54034 => x"082082",
   54035 => x"082041",
   54036 => x"041041",
   54037 => x"041041",
   54038 => x"041041",
   54039 => x"041041",
   54040 => x"041041",
   54041 => x"041041",
   54042 => x"041041",
   54043 => x"041041",
   54044 => x"041041",
   54045 => x"041041",
   54046 => x"041041",
   54047 => x"041041",
   54048 => x"041041",
   54049 => x"041041",
   54050 => x"041041",
   54051 => x"041041",
   54052 => x"041041",
   54053 => x"041041",
   54054 => x"041041",
   54055 => x"041041",
   54056 => x"041041",
   54057 => x"041041",
   54058 => x"041000",
   54059 => x"000000",
   54060 => x"000000",
   54061 => x"000000",
   54062 => x"000000",
   54063 => x"000000",
   54064 => x"000000",
   54065 => x"000000",
   54066 => x"000000",
   54067 => x"000000",
   54068 => x"000000",
   54069 => x"00057f",
   54070 => x"ffffff",
   54071 => x"ffffff",
   54072 => x"ffffff",
   54073 => x"ffffd5",
   54074 => x"00002a",
   54075 => x"ffffff",
   54076 => x"ffffff",
   54077 => x"fea540",
   54078 => x"00056a",
   54079 => x"ffffff",
   54080 => x"ffffff",
   54081 => x"ffffff",
   54082 => x"ffffff",
   54083 => x"ffffff",
   54084 => x"ffffff",
   54085 => x"ffffff",
   54086 => x"ffffff",
   54087 => x"ffffff",
   54088 => x"ffffff",
   54089 => x"ffffff",
   54090 => x"ffffff",
   54091 => x"ffffff",
   54092 => x"ffffff",
   54093 => x"ffffff",
   54094 => x"ffffff",
   54095 => x"ffffff",
   54096 => x"ffffff",
   54097 => x"ffffff",
   54098 => x"ffffff",
   54099 => x"ffffff",
   54100 => x"ffffff",
   54101 => x"ffffff",
   54102 => x"ffffff",
   54103 => x"ffffff",
   54104 => x"ffffff",
   54105 => x"ffffff",
   54106 => x"ffffff",
   54107 => x"ffffff",
   54108 => x"ffffff",
   54109 => x"ffffff",
   54110 => x"ffffff",
   54111 => x"ffffff",
   54112 => x"ffffff",
   54113 => x"ffffff",
   54114 => x"ffffff",
   54115 => x"ffffff",
   54116 => x"ffffff",
   54117 => x"ffffff",
   54118 => x"ffffff",
   54119 => x"ffffff",
   54120 => x"ffffff",
   54121 => x"ffffff",
   54122 => x"ffffff",
   54123 => x"ffffff",
   54124 => x"ffffff",
   54125 => x"ffffff",
   54126 => x"ffffff",
   54127 => x"ffffff",
   54128 => x"ffffff",
   54129 => x"ffffff",
   54130 => x"ffffff",
   54131 => x"ffffff",
   54132 => x"ffffff",
   54133 => x"ffffff",
   54134 => x"ffffff",
   54135 => x"ffffff",
   54136 => x"ffffff",
   54137 => x"ffffff",
   54138 => x"ffffff",
   54139 => x"ffffff",
   54140 => x"ffffff",
   54141 => x"ffffff",
   54142 => x"ffffff",
   54143 => x"ffffff",
   54144 => x"ffffff",
   54145 => x"ffffff",
   54146 => x"ffffff",
   54147 => x"ffffff",
   54148 => x"ffffff",
   54149 => x"fffa95",
   54150 => x"abffff",
   54151 => x"ffffff",
   54152 => x"ffffff",
   54153 => x"ffffff",
   54154 => x"ffffff",
   54155 => x"ffffff",
   54156 => x"ffffff",
   54157 => x"ffffff",
   54158 => x"ffffff",
   54159 => x"ffffff",
   54160 => x"ffffff",
   54161 => x"fffac3",
   54162 => x"0c30c3",
   54163 => x"0c30c3",
   54164 => x"0c30c3",
   54165 => x"0c30c3",
   54166 => x"0c30c3",
   54167 => x"0c30c3",
   54168 => x"0c30c3",
   54169 => x"0c30c3",
   54170 => x"0c30c3",
   54171 => x"0c30c3",
   54172 => x"0c30c3",
   54173 => x"082082",
   54174 => x"082082",
   54175 => x"082082",
   54176 => x"082082",
   54177 => x"082082",
   54178 => x"082082",
   54179 => x"082082",
   54180 => x"082082",
   54181 => x"082082",
   54182 => x"082082",
   54183 => x"082082",
   54184 => x"082082",
   54185 => x"082082",
   54186 => x"082082",
   54187 => x"082082",
   54188 => x"082082",
   54189 => x"082082",
   54190 => x"082082",
   54191 => x"082082",
   54192 => x"082082",
   54193 => x"082082",
   54194 => x"082082",
   54195 => x"082041",
   54196 => x"041041",
   54197 => x"041041",
   54198 => x"041041",
   54199 => x"041041",
   54200 => x"041041",
   54201 => x"041041",
   54202 => x"041041",
   54203 => x"041041",
   54204 => x"041041",
   54205 => x"041041",
   54206 => x"041041",
   54207 => x"041041",
   54208 => x"041041",
   54209 => x"041041",
   54210 => x"041041",
   54211 => x"041041",
   54212 => x"041041",
   54213 => x"041041",
   54214 => x"041041",
   54215 => x"041041",
   54216 => x"041041",
   54217 => x"041041",
   54218 => x"041000",
   54219 => x"000000",
   54220 => x"000000",
   54221 => x"000000",
   54222 => x"000000",
   54223 => x"000000",
   54224 => x"000000",
   54225 => x"000000",
   54226 => x"000000",
   54227 => x"000000",
   54228 => x"000000",
   54229 => x"00057f",
   54230 => x"ffffff",
   54231 => x"ffffff",
   54232 => x"ffffff",
   54233 => x"ffffd5",
   54234 => x"00002a",
   54235 => x"ffffff",
   54236 => x"ffffff",
   54237 => x"ffffd5",
   54238 => x"000015",
   54239 => x"ffffff",
   54240 => x"ffffff",
   54241 => x"ffffff",
   54242 => x"ffffff",
   54243 => x"ffffff",
   54244 => x"ffffff",
   54245 => x"ffffff",
   54246 => x"ffffff",
   54247 => x"ffffff",
   54248 => x"ffffff",
   54249 => x"ffffff",
   54250 => x"ffffff",
   54251 => x"ffffff",
   54252 => x"ffffff",
   54253 => x"ffffff",
   54254 => x"ffffff",
   54255 => x"ffffff",
   54256 => x"ffffff",
   54257 => x"ffffff",
   54258 => x"ffffff",
   54259 => x"ffffff",
   54260 => x"ffffff",
   54261 => x"ffffff",
   54262 => x"ffffff",
   54263 => x"ffffff",
   54264 => x"ffffff",
   54265 => x"ffffff",
   54266 => x"ffffff",
   54267 => x"ffffff",
   54268 => x"ffffff",
   54269 => x"ffffff",
   54270 => x"ffffff",
   54271 => x"ffffff",
   54272 => x"ffffff",
   54273 => x"ffffff",
   54274 => x"ffffff",
   54275 => x"ffffff",
   54276 => x"ffffff",
   54277 => x"ffffff",
   54278 => x"ffffff",
   54279 => x"ffffff",
   54280 => x"ffffff",
   54281 => x"ffffff",
   54282 => x"ffffff",
   54283 => x"ffffff",
   54284 => x"ffffff",
   54285 => x"ffffff",
   54286 => x"ffffff",
   54287 => x"ffffff",
   54288 => x"ffffff",
   54289 => x"ffffff",
   54290 => x"ffffff",
   54291 => x"ffffff",
   54292 => x"ffffff",
   54293 => x"ffffff",
   54294 => x"ffffff",
   54295 => x"ffffff",
   54296 => x"ffffff",
   54297 => x"ffffff",
   54298 => x"ffffff",
   54299 => x"ffffff",
   54300 => x"ffffff",
   54301 => x"ffffff",
   54302 => x"ffffff",
   54303 => x"ffffff",
   54304 => x"ffffff",
   54305 => x"ffffff",
   54306 => x"ffffff",
   54307 => x"ffffff",
   54308 => x"ffffff",
   54309 => x"fffa95",
   54310 => x"abffff",
   54311 => x"ffffff",
   54312 => x"ffffff",
   54313 => x"ffffff",
   54314 => x"ffffff",
   54315 => x"ffffff",
   54316 => x"ffffff",
   54317 => x"ffffff",
   54318 => x"ffffff",
   54319 => x"ffffff",
   54320 => x"ffffff",
   54321 => x"fffac3",
   54322 => x"0c30c3",
   54323 => x"0c30c3",
   54324 => x"0c30c3",
   54325 => x"0c30c3",
   54326 => x"0c30c3",
   54327 => x"0c30c3",
   54328 => x"0c30c3",
   54329 => x"0c30c3",
   54330 => x"0c30c3",
   54331 => x"0c30c3",
   54332 => x"0c30c3",
   54333 => x"082082",
   54334 => x"082082",
   54335 => x"082082",
   54336 => x"082082",
   54337 => x"082082",
   54338 => x"082082",
   54339 => x"082082",
   54340 => x"082082",
   54341 => x"082082",
   54342 => x"082082",
   54343 => x"082082",
   54344 => x"082082",
   54345 => x"082082",
   54346 => x"082082",
   54347 => x"082082",
   54348 => x"082082",
   54349 => x"082082",
   54350 => x"082082",
   54351 => x"082082",
   54352 => x"082082",
   54353 => x"082082",
   54354 => x"082082",
   54355 => x"082041",
   54356 => x"041041",
   54357 => x"041041",
   54358 => x"041041",
   54359 => x"041041",
   54360 => x"041041",
   54361 => x"041041",
   54362 => x"041041",
   54363 => x"041041",
   54364 => x"041041",
   54365 => x"041041",
   54366 => x"041041",
   54367 => x"041041",
   54368 => x"041041",
   54369 => x"041041",
   54370 => x"041041",
   54371 => x"041041",
   54372 => x"041041",
   54373 => x"041041",
   54374 => x"041041",
   54375 => x"041041",
   54376 => x"041041",
   54377 => x"041041",
   54378 => x"041000",
   54379 => x"000000",
   54380 => x"000000",
   54381 => x"000000",
   54382 => x"000000",
   54383 => x"000000",
   54384 => x"000000",
   54385 => x"000000",
   54386 => x"000000",
   54387 => x"000000",
   54388 => x"000000",
   54389 => x"00057f",
   54390 => x"ffffff",
   54391 => x"ffffff",
   54392 => x"ffffff",
   54393 => x"ffffd5",
   54394 => x"00002a",
   54395 => x"ffffff",
   54396 => x"ffffff",
   54397 => x"ffffea",
   54398 => x"000000",
   54399 => x"abffff",
   54400 => x"ffffff",
   54401 => x"ffffff",
   54402 => x"ffffff",
   54403 => x"ffffff",
   54404 => x"ffffff",
   54405 => x"ffffff",
   54406 => x"ffffff",
   54407 => x"ffffff",
   54408 => x"ffffff",
   54409 => x"ffffff",
   54410 => x"ffffff",
   54411 => x"ffffff",
   54412 => x"ffffff",
   54413 => x"ffffff",
   54414 => x"ffffff",
   54415 => x"ffffff",
   54416 => x"ffffff",
   54417 => x"ffffff",
   54418 => x"ffffff",
   54419 => x"ffffff",
   54420 => x"ffffff",
   54421 => x"ffffff",
   54422 => x"ffffff",
   54423 => x"ffffff",
   54424 => x"ffffff",
   54425 => x"ffffff",
   54426 => x"ffffff",
   54427 => x"ffffff",
   54428 => x"ffffff",
   54429 => x"ffffff",
   54430 => x"ffffff",
   54431 => x"ffffff",
   54432 => x"ffffff",
   54433 => x"ffffff",
   54434 => x"ffffff",
   54435 => x"ffffff",
   54436 => x"ffffff",
   54437 => x"ffffff",
   54438 => x"ffffff",
   54439 => x"ffffff",
   54440 => x"ffffff",
   54441 => x"ffffff",
   54442 => x"ffffff",
   54443 => x"ffffff",
   54444 => x"ffffff",
   54445 => x"ffffff",
   54446 => x"ffffff",
   54447 => x"ffffff",
   54448 => x"ffffff",
   54449 => x"ffffff",
   54450 => x"ffffff",
   54451 => x"ffffff",
   54452 => x"ffffff",
   54453 => x"ffffff",
   54454 => x"ffffff",
   54455 => x"ffffff",
   54456 => x"ffffff",
   54457 => x"ffffff",
   54458 => x"ffffff",
   54459 => x"ffffff",
   54460 => x"ffffff",
   54461 => x"ffffff",
   54462 => x"ffffff",
   54463 => x"ffffff",
   54464 => x"ffffff",
   54465 => x"ffffff",
   54466 => x"ffffff",
   54467 => x"ffffff",
   54468 => x"ffffff",
   54469 => x"fffa95",
   54470 => x"abffff",
   54471 => x"ffffff",
   54472 => x"ffffff",
   54473 => x"ffffff",
   54474 => x"ffffff",
   54475 => x"ffffff",
   54476 => x"ffffff",
   54477 => x"ffffff",
   54478 => x"ffffff",
   54479 => x"ffffff",
   54480 => x"ffffff",
   54481 => x"fffac3",
   54482 => x"0c30c3",
   54483 => x"0c30c3",
   54484 => x"0c30c3",
   54485 => x"0c30c3",
   54486 => x"0c30c3",
   54487 => x"0c30c3",
   54488 => x"0c30c3",
   54489 => x"0c30c3",
   54490 => x"0c30c3",
   54491 => x"0c30c3",
   54492 => x"0c30c3",
   54493 => x"082082",
   54494 => x"082082",
   54495 => x"082082",
   54496 => x"082082",
   54497 => x"082082",
   54498 => x"082082",
   54499 => x"082082",
   54500 => x"082082",
   54501 => x"082082",
   54502 => x"082082",
   54503 => x"082082",
   54504 => x"082082",
   54505 => x"082082",
   54506 => x"082082",
   54507 => x"082082",
   54508 => x"082082",
   54509 => x"082082",
   54510 => x"082082",
   54511 => x"082082",
   54512 => x"082082",
   54513 => x"082082",
   54514 => x"082082",
   54515 => x"082041",
   54516 => x"041041",
   54517 => x"041041",
   54518 => x"041041",
   54519 => x"041041",
   54520 => x"041041",
   54521 => x"041041",
   54522 => x"041041",
   54523 => x"041041",
   54524 => x"041041",
   54525 => x"041041",
   54526 => x"041041",
   54527 => x"041041",
   54528 => x"041041",
   54529 => x"041041",
   54530 => x"041041",
   54531 => x"041041",
   54532 => x"041041",
   54533 => x"041041",
   54534 => x"041041",
   54535 => x"041041",
   54536 => x"041041",
   54537 => x"041041",
   54538 => x"041000",
   54539 => x"000000",
   54540 => x"000000",
   54541 => x"000000",
   54542 => x"000000",
   54543 => x"000000",
   54544 => x"000000",
   54545 => x"000000",
   54546 => x"000000",
   54547 => x"000000",
   54548 => x"000000",
   54549 => x"00057f",
   54550 => x"ffffff",
   54551 => x"ffffff",
   54552 => x"ffffff",
   54553 => x"ffffd5",
   54554 => x"00002a",
   54555 => x"ffffff",
   54556 => x"ffffff",
   54557 => x"ffffff",
   54558 => x"540000",
   54559 => x"57ffff",
   54560 => x"ffffff",
   54561 => x"ffffff",
   54562 => x"ffffff",
   54563 => x"ffffff",
   54564 => x"ffffff",
   54565 => x"ffffff",
   54566 => x"ffffff",
   54567 => x"ffffff",
   54568 => x"ffffff",
   54569 => x"ffffff",
   54570 => x"ffffff",
   54571 => x"ffffff",
   54572 => x"ffffff",
   54573 => x"ffffff",
   54574 => x"ffffff",
   54575 => x"ffffff",
   54576 => x"ffffff",
   54577 => x"ffffff",
   54578 => x"ffffff",
   54579 => x"ffffff",
   54580 => x"ffffff",
   54581 => x"ffffff",
   54582 => x"ffffff",
   54583 => x"ffffff",
   54584 => x"ffffff",
   54585 => x"ffffff",
   54586 => x"ffffff",
   54587 => x"ffffff",
   54588 => x"ffffff",
   54589 => x"ffffff",
   54590 => x"ffffff",
   54591 => x"ffffff",
   54592 => x"ffffff",
   54593 => x"ffffff",
   54594 => x"ffffff",
   54595 => x"ffffff",
   54596 => x"ffffff",
   54597 => x"ffffff",
   54598 => x"ffffff",
   54599 => x"ffffff",
   54600 => x"ffffff",
   54601 => x"ffffff",
   54602 => x"ffffff",
   54603 => x"ffffff",
   54604 => x"ffffff",
   54605 => x"ffffff",
   54606 => x"ffffff",
   54607 => x"ffffff",
   54608 => x"ffffff",
   54609 => x"ffffff",
   54610 => x"ffffff",
   54611 => x"ffffff",
   54612 => x"ffffff",
   54613 => x"ffffff",
   54614 => x"ffffff",
   54615 => x"ffffff",
   54616 => x"ffffff",
   54617 => x"ffffff",
   54618 => x"ffffff",
   54619 => x"ffffff",
   54620 => x"ffffff",
   54621 => x"ffffff",
   54622 => x"ffffff",
   54623 => x"ffffff",
   54624 => x"ffffff",
   54625 => x"ffffff",
   54626 => x"ffffff",
   54627 => x"ffffff",
   54628 => x"ffffff",
   54629 => x"fffa95",
   54630 => x"abffff",
   54631 => x"ffffff",
   54632 => x"ffffff",
   54633 => x"ffffff",
   54634 => x"ffffff",
   54635 => x"ffffff",
   54636 => x"ffffff",
   54637 => x"ffffff",
   54638 => x"ffffff",
   54639 => x"ffffff",
   54640 => x"ffffff",
   54641 => x"fffac3",
   54642 => x"0c30c3",
   54643 => x"0c30c3",
   54644 => x"0c30c3",
   54645 => x"0c30c3",
   54646 => x"0c30c3",
   54647 => x"0c30c3",
   54648 => x"0c30c3",
   54649 => x"0c30c3",
   54650 => x"0c30c3",
   54651 => x"0c30c3",
   54652 => x"0c30c3",
   54653 => x"082082",
   54654 => x"082082",
   54655 => x"082082",
   54656 => x"082082",
   54657 => x"082082",
   54658 => x"082082",
   54659 => x"082082",
   54660 => x"082082",
   54661 => x"082082",
   54662 => x"082082",
   54663 => x"082082",
   54664 => x"082082",
   54665 => x"082082",
   54666 => x"082082",
   54667 => x"082082",
   54668 => x"082082",
   54669 => x"082082",
   54670 => x"082082",
   54671 => x"082082",
   54672 => x"082082",
   54673 => x"082082",
   54674 => x"082082",
   54675 => x"082041",
   54676 => x"041041",
   54677 => x"041041",
   54678 => x"041041",
   54679 => x"041041",
   54680 => x"041041",
   54681 => x"041041",
   54682 => x"041041",
   54683 => x"041041",
   54684 => x"041041",
   54685 => x"041041",
   54686 => x"041041",
   54687 => x"041041",
   54688 => x"041041",
   54689 => x"041041",
   54690 => x"041041",
   54691 => x"041041",
   54692 => x"041041",
   54693 => x"041041",
   54694 => x"041041",
   54695 => x"041041",
   54696 => x"041041",
   54697 => x"041041",
   54698 => x"041000",
   54699 => x"000000",
   54700 => x"000000",
   54701 => x"000000",
   54702 => x"000000",
   54703 => x"000000",
   54704 => x"000000",
   54705 => x"000000",
   54706 => x"000000",
   54707 => x"000000",
   54708 => x"000000",
   54709 => x"00057f",
   54710 => x"ffffff",
   54711 => x"ffffff",
   54712 => x"ffffff",
   54713 => x"ffffd5",
   54714 => x"00002a",
   54715 => x"ffffff",
   54716 => x"ffffff",
   54717 => x"ffffff",
   54718 => x"540000",
   54719 => x"57ffff",
   54720 => x"ffffff",
   54721 => x"ffffff",
   54722 => x"ffffff",
   54723 => x"ffffff",
   54724 => x"ffffff",
   54725 => x"ffffff",
   54726 => x"ffffff",
   54727 => x"ffffff",
   54728 => x"ffffff",
   54729 => x"ffffff",
   54730 => x"ffffff",
   54731 => x"ffffff",
   54732 => x"ffffff",
   54733 => x"ffffff",
   54734 => x"ffffff",
   54735 => x"ffffff",
   54736 => x"ffffff",
   54737 => x"ffffff",
   54738 => x"ffffff",
   54739 => x"ffffff",
   54740 => x"ffffff",
   54741 => x"ffffff",
   54742 => x"ffffff",
   54743 => x"ffffff",
   54744 => x"ffffff",
   54745 => x"ffffff",
   54746 => x"ffffff",
   54747 => x"ffffff",
   54748 => x"ffffff",
   54749 => x"ffffff",
   54750 => x"ffffff",
   54751 => x"ffffff",
   54752 => x"ffffff",
   54753 => x"ffffff",
   54754 => x"ffffff",
   54755 => x"ffffff",
   54756 => x"ffffff",
   54757 => x"ffffff",
   54758 => x"ffffff",
   54759 => x"ffffff",
   54760 => x"ffffff",
   54761 => x"ffffff",
   54762 => x"ffffff",
   54763 => x"ffffff",
   54764 => x"ffffff",
   54765 => x"ffffff",
   54766 => x"ffffff",
   54767 => x"ffffff",
   54768 => x"ffffff",
   54769 => x"ffffff",
   54770 => x"ffffff",
   54771 => x"ffffff",
   54772 => x"ffffff",
   54773 => x"ffffff",
   54774 => x"ffffff",
   54775 => x"ffffff",
   54776 => x"ffffff",
   54777 => x"ffffff",
   54778 => x"ffffff",
   54779 => x"ffffff",
   54780 => x"ffffff",
   54781 => x"ffffff",
   54782 => x"ffffff",
   54783 => x"ffffff",
   54784 => x"ffffff",
   54785 => x"ffffff",
   54786 => x"ffffff",
   54787 => x"ffffff",
   54788 => x"ffffff",
   54789 => x"fffa95",
   54790 => x"abffff",
   54791 => x"ffffff",
   54792 => x"ffffff",
   54793 => x"ffffff",
   54794 => x"ffffff",
   54795 => x"ffffff",
   54796 => x"ffffff",
   54797 => x"ffffff",
   54798 => x"ffffff",
   54799 => x"ffffff",
   54800 => x"ffffff",
   54801 => x"fffac3",
   54802 => x"0c30c3",
   54803 => x"0c30c3",
   54804 => x"0c30c3",
   54805 => x"0c30c3",
   54806 => x"0c30c3",
   54807 => x"0c30c3",
   54808 => x"0c30c3",
   54809 => x"0c30c3",
   54810 => x"0c30c3",
   54811 => x"0c30c3",
   54812 => x"0c30c3",
   54813 => x"082082",
   54814 => x"082082",
   54815 => x"082082",
   54816 => x"082082",
   54817 => x"082082",
   54818 => x"082082",
   54819 => x"082082",
   54820 => x"082082",
   54821 => x"082082",
   54822 => x"082082",
   54823 => x"082082",
   54824 => x"082082",
   54825 => x"082082",
   54826 => x"082082",
   54827 => x"082082",
   54828 => x"082082",
   54829 => x"082082",
   54830 => x"082082",
   54831 => x"082082",
   54832 => x"082082",
   54833 => x"082082",
   54834 => x"082082",
   54835 => x"082041",
   54836 => x"041041",
   54837 => x"041041",
   54838 => x"041041",
   54839 => x"041041",
   54840 => x"041041",
   54841 => x"041041",
   54842 => x"041041",
   54843 => x"041041",
   54844 => x"041041",
   54845 => x"041041",
   54846 => x"041041",
   54847 => x"041041",
   54848 => x"041041",
   54849 => x"041041",
   54850 => x"041041",
   54851 => x"041041",
   54852 => x"041041",
   54853 => x"041041",
   54854 => x"041041",
   54855 => x"041041",
   54856 => x"041041",
   54857 => x"041041",
   54858 => x"041000",
   54859 => x"000000",
   54860 => x"000000",
   54861 => x"000000",
   54862 => x"000000",
   54863 => x"000000",
   54864 => x"000000",
   54865 => x"000000",
   54866 => x"000000",
   54867 => x"000000",
   54868 => x"000000",
   54869 => x"00057f",
   54870 => x"ffffff",
   54871 => x"ffffff",
   54872 => x"ffffff",
   54873 => x"ffffd5",
   54874 => x"00002a",
   54875 => x"ffffff",
   54876 => x"ffffff",
   54877 => x"ffffff",
   54878 => x"540000",
   54879 => x"57ffff",
   54880 => x"ffffff",
   54881 => x"ffffff",
   54882 => x"ffffff",
   54883 => x"ffffff",
   54884 => x"ffffff",
   54885 => x"ffffff",
   54886 => x"ffffff",
   54887 => x"ffffff",
   54888 => x"ffffff",
   54889 => x"ffffff",
   54890 => x"ffffff",
   54891 => x"ffffff",
   54892 => x"ffffff",
   54893 => x"ffffff",
   54894 => x"ffffff",
   54895 => x"ffffff",
   54896 => x"ffffff",
   54897 => x"ffffff",
   54898 => x"ffffff",
   54899 => x"ffffff",
   54900 => x"ffffff",
   54901 => x"ffffff",
   54902 => x"ffffff",
   54903 => x"ffffff",
   54904 => x"ffffff",
   54905 => x"ffffff",
   54906 => x"ffffff",
   54907 => x"ffffff",
   54908 => x"ffffff",
   54909 => x"ffffff",
   54910 => x"ffffff",
   54911 => x"ffffff",
   54912 => x"ffffff",
   54913 => x"ffffff",
   54914 => x"ffffff",
   54915 => x"ffffff",
   54916 => x"ffffff",
   54917 => x"ffffff",
   54918 => x"ffffff",
   54919 => x"ffffff",
   54920 => x"ffffff",
   54921 => x"ffffff",
   54922 => x"ffffff",
   54923 => x"ffffff",
   54924 => x"ffffff",
   54925 => x"ffffff",
   54926 => x"ffffff",
   54927 => x"ffffff",
   54928 => x"ffffff",
   54929 => x"ffffff",
   54930 => x"ffffff",
   54931 => x"ffffff",
   54932 => x"ffffff",
   54933 => x"ffffff",
   54934 => x"ffffff",
   54935 => x"ffffff",
   54936 => x"ffffff",
   54937 => x"ffffff",
   54938 => x"ffffff",
   54939 => x"ffffff",
   54940 => x"ffffff",
   54941 => x"ffffff",
   54942 => x"ffffff",
   54943 => x"ffffff",
   54944 => x"ffffff",
   54945 => x"ffffff",
   54946 => x"ffffff",
   54947 => x"ffffff",
   54948 => x"ffffff",
   54949 => x"fffa95",
   54950 => x"abffff",
   54951 => x"ffffff",
   54952 => x"ffffff",
   54953 => x"ffffff",
   54954 => x"ffffff",
   54955 => x"ffffff",
   54956 => x"ffffff",
   54957 => x"ffffff",
   54958 => x"ffffff",
   54959 => x"ffffff",
   54960 => x"ffffff",
   54961 => x"fffac3",
   54962 => x"0c30c3",
   54963 => x"0c30c3",
   54964 => x"0c30c3",
   54965 => x"0c30c3",
   54966 => x"0c30c3",
   54967 => x"0c30c3",
   54968 => x"0c30c3",
   54969 => x"0c30c3",
   54970 => x"0c30c3",
   54971 => x"0c30c3",
   54972 => x"0c30c3",
   54973 => x"082082",
   54974 => x"082082",
   54975 => x"082082",
   54976 => x"082082",
   54977 => x"082082",
   54978 => x"082082",
   54979 => x"082082",
   54980 => x"082082",
   54981 => x"082082",
   54982 => x"082082",
   54983 => x"082082",
   54984 => x"082082",
   54985 => x"082082",
   54986 => x"082082",
   54987 => x"082082",
   54988 => x"082082",
   54989 => x"082082",
   54990 => x"082082",
   54991 => x"082082",
   54992 => x"082082",
   54993 => x"082082",
   54994 => x"082082",
   54995 => x"082041",
   54996 => x"041041",
   54997 => x"041041",
   54998 => x"041041",
   54999 => x"041041",
   55000 => x"041041",
   55001 => x"041041",
   55002 => x"041041",
   55003 => x"041041",
   55004 => x"041041",
   55005 => x"041041",
   55006 => x"041041",
   55007 => x"041041",
   55008 => x"041041",
   55009 => x"041041",
   55010 => x"041041",
   55011 => x"041041",
   55012 => x"041041",
   55013 => x"041041",
   55014 => x"041041",
   55015 => x"041041",
   55016 => x"041041",
   55017 => x"041041",
   55018 => x"041000",
   55019 => x"000000",
   55020 => x"000000",
   55021 => x"000000",
   55022 => x"000000",
   55023 => x"000000",
   55024 => x"000000",
   55025 => x"000000",
   55026 => x"000000",
   55027 => x"000000",
   55028 => x"000000",
   55029 => x"00057f",
   55030 => x"ffffff",
   55031 => x"ffffff",
   55032 => x"ffffff",
   55033 => x"ffffd5",
   55034 => x"00002a",
   55035 => x"ffffff",
   55036 => x"ffffff",
   55037 => x"ffffff",
   55038 => x"540000",
   55039 => x"57ffff",
   55040 => x"ffffff",
   55041 => x"ffffff",
   55042 => x"ffffff",
   55043 => x"ffffff",
   55044 => x"ffffff",
   55045 => x"ffffff",
   55046 => x"ffffff",
   55047 => x"ffffff",
   55048 => x"ffffff",
   55049 => x"ffffff",
   55050 => x"ffffff",
   55051 => x"ffffff",
   55052 => x"ffffff",
   55053 => x"ffffff",
   55054 => x"ffffff",
   55055 => x"ffffff",
   55056 => x"ffffff",
   55057 => x"ffffff",
   55058 => x"ffffff",
   55059 => x"ffffff",
   55060 => x"ffffff",
   55061 => x"ffffff",
   55062 => x"ffffff",
   55063 => x"ffffff",
   55064 => x"ffffff",
   55065 => x"ffffff",
   55066 => x"ffffff",
   55067 => x"ffffff",
   55068 => x"ffffff",
   55069 => x"ffffff",
   55070 => x"ffffff",
   55071 => x"ffffff",
   55072 => x"ffffff",
   55073 => x"ffffff",
   55074 => x"ffffff",
   55075 => x"ffffff",
   55076 => x"ffffff",
   55077 => x"ffffff",
   55078 => x"ffffff",
   55079 => x"ffffff",
   55080 => x"ffffff",
   55081 => x"ffffff",
   55082 => x"ffffff",
   55083 => x"ffffff",
   55084 => x"ffffff",
   55085 => x"ffffff",
   55086 => x"ffffff",
   55087 => x"ffffff",
   55088 => x"ffffff",
   55089 => x"ffffff",
   55090 => x"ffffff",
   55091 => x"ffffff",
   55092 => x"ffffff",
   55093 => x"ffffff",
   55094 => x"ffffff",
   55095 => x"ffffff",
   55096 => x"ffffff",
   55097 => x"ffffff",
   55098 => x"ffffff",
   55099 => x"ffffff",
   55100 => x"ffffff",
   55101 => x"ffffff",
   55102 => x"ffffff",
   55103 => x"ffffff",
   55104 => x"ffffff",
   55105 => x"ffffff",
   55106 => x"ffffff",
   55107 => x"ffffff",
   55108 => x"ffffff",
   55109 => x"fffa95",
   55110 => x"abffff",
   55111 => x"ffffff",
   55112 => x"ffffff",
   55113 => x"ffffff",
   55114 => x"ffffff",
   55115 => x"ffffff",
   55116 => x"ffffff",
   55117 => x"ffffff",
   55118 => x"ffffff",
   55119 => x"ffffff",
   55120 => x"ffffff",
   55121 => x"fffac3",
   55122 => x"0c30c3",
   55123 => x"0c30c3",
   55124 => x"0c30c3",
   55125 => x"0c30c3",
   55126 => x"0c30c3",
   55127 => x"0c30c3",
   55128 => x"0c30c3",
   55129 => x"0c30c3",
   55130 => x"0c30c3",
   55131 => x"0c30c3",
   55132 => x"0c30c3",
   55133 => x"082082",
   55134 => x"082082",
   55135 => x"082082",
   55136 => x"082082",
   55137 => x"082082",
   55138 => x"082082",
   55139 => x"082082",
   55140 => x"082082",
   55141 => x"082082",
   55142 => x"082082",
   55143 => x"082082",
   55144 => x"082082",
   55145 => x"082082",
   55146 => x"082082",
   55147 => x"082082",
   55148 => x"082082",
   55149 => x"082082",
   55150 => x"082082",
   55151 => x"082082",
   55152 => x"082082",
   55153 => x"082082",
   55154 => x"082082",
   55155 => x"082041",
   55156 => x"041041",
   55157 => x"041041",
   55158 => x"041041",
   55159 => x"041041",
   55160 => x"041041",
   55161 => x"041041",
   55162 => x"041041",
   55163 => x"041041",
   55164 => x"041041",
   55165 => x"041041",
   55166 => x"041041",
   55167 => x"041041",
   55168 => x"041041",
   55169 => x"041041",
   55170 => x"041041",
   55171 => x"041041",
   55172 => x"041041",
   55173 => x"041041",
   55174 => x"041041",
   55175 => x"041041",
   55176 => x"041041",
   55177 => x"041041",
   55178 => x"041000",
   55179 => x"000000",
   55180 => x"000000",
   55181 => x"000000",
   55182 => x"000000",
   55183 => x"000000",
   55184 => x"000000",
   55185 => x"000000",
   55186 => x"000000",
   55187 => x"000000",
   55188 => x"000000",
   55189 => x"00057f",
   55190 => x"ffffff",
   55191 => x"ffffff",
   55192 => x"ffffff",
   55193 => x"ffffd5",
   55194 => x"00002a",
   55195 => x"ffffff",
   55196 => x"ffffff",
   55197 => x"ffffea",
   55198 => x"540000",
   55199 => x"57ffff",
   55200 => x"ffffff",
   55201 => x"ffffff",
   55202 => x"ffffff",
   55203 => x"ffffff",
   55204 => x"ffffff",
   55205 => x"ffffff",
   55206 => x"ffffff",
   55207 => x"ffffff",
   55208 => x"ffffff",
   55209 => x"ffffff",
   55210 => x"ffffff",
   55211 => x"ffffff",
   55212 => x"ffffff",
   55213 => x"ffffff",
   55214 => x"ffffff",
   55215 => x"ffffff",
   55216 => x"ffffff",
   55217 => x"ffffff",
   55218 => x"ffffff",
   55219 => x"ffffff",
   55220 => x"ffffff",
   55221 => x"ffffff",
   55222 => x"ffffff",
   55223 => x"ffffff",
   55224 => x"ffffff",
   55225 => x"ffffff",
   55226 => x"ffffff",
   55227 => x"ffffff",
   55228 => x"ffffff",
   55229 => x"ffffff",
   55230 => x"ffffff",
   55231 => x"ffffff",
   55232 => x"ffffff",
   55233 => x"ffffff",
   55234 => x"ffffff",
   55235 => x"ffffff",
   55236 => x"ffffff",
   55237 => x"ffffff",
   55238 => x"ffffff",
   55239 => x"ffffff",
   55240 => x"ffffff",
   55241 => x"ffffff",
   55242 => x"ffffff",
   55243 => x"ffffff",
   55244 => x"ffffff",
   55245 => x"ffffff",
   55246 => x"ffffff",
   55247 => x"ffffff",
   55248 => x"ffffff",
   55249 => x"ffffff",
   55250 => x"ffffff",
   55251 => x"ffffff",
   55252 => x"ffffff",
   55253 => x"ffffff",
   55254 => x"ffffff",
   55255 => x"ffffff",
   55256 => x"ffffff",
   55257 => x"ffffff",
   55258 => x"ffffff",
   55259 => x"ffffff",
   55260 => x"ffffff",
   55261 => x"ffffff",
   55262 => x"ffffff",
   55263 => x"ffffff",
   55264 => x"ffffff",
   55265 => x"ffffff",
   55266 => x"ffffff",
   55267 => x"ffffff",
   55268 => x"ffffff",
   55269 => x"fffa95",
   55270 => x"abffff",
   55271 => x"ffffff",
   55272 => x"ffffff",
   55273 => x"ffffff",
   55274 => x"ffffff",
   55275 => x"ffffff",
   55276 => x"ffffff",
   55277 => x"ffffff",
   55278 => x"ffffff",
   55279 => x"ffffff",
   55280 => x"ffffff",
   55281 => x"fffac3",
   55282 => x"0c30c3",
   55283 => x"0c30c3",
   55284 => x"0c30c3",
   55285 => x"0c30c3",
   55286 => x"0c30c3",
   55287 => x"0c30c3",
   55288 => x"0c30c3",
   55289 => x"0c30c3",
   55290 => x"0c30c3",
   55291 => x"0c30c3",
   55292 => x"0c30c3",
   55293 => x"082082",
   55294 => x"082082",
   55295 => x"082082",
   55296 => x"082082",
   55297 => x"082082",
   55298 => x"082082",
   55299 => x"082082",
   55300 => x"082082",
   55301 => x"082082",
   55302 => x"082082",
   55303 => x"082082",
   55304 => x"082082",
   55305 => x"082082",
   55306 => x"082082",
   55307 => x"082082",
   55308 => x"082082",
   55309 => x"082082",
   55310 => x"082082",
   55311 => x"082082",
   55312 => x"082082",
   55313 => x"082082",
   55314 => x"082082",
   55315 => x"082041",
   55316 => x"041041",
   55317 => x"041041",
   55318 => x"041041",
   55319 => x"041041",
   55320 => x"041041",
   55321 => x"041041",
   55322 => x"041041",
   55323 => x"041041",
   55324 => x"041041",
   55325 => x"041041",
   55326 => x"041041",
   55327 => x"041041",
   55328 => x"041041",
   55329 => x"041041",
   55330 => x"041041",
   55331 => x"041041",
   55332 => x"041041",
   55333 => x"041041",
   55334 => x"041041",
   55335 => x"041041",
   55336 => x"041041",
   55337 => x"041041",
   55338 => x"041000",
   55339 => x"000000",
   55340 => x"000000",
   55341 => x"000000",
   55342 => x"000000",
   55343 => x"000000",
   55344 => x"000000",
   55345 => x"000000",
   55346 => x"000000",
   55347 => x"000000",
   55348 => x"000000",
   55349 => x"00057f",
   55350 => x"ffffff",
   55351 => x"ffffff",
   55352 => x"ffffff",
   55353 => x"ffffd5",
   55354 => x"00002a",
   55355 => x"ffffff",
   55356 => x"ffffff",
   55357 => x"ffffd5",
   55358 => x"000000",
   55359 => x"abffff",
   55360 => x"ffffff",
   55361 => x"ffffff",
   55362 => x"ffffff",
   55363 => x"ffffff",
   55364 => x"ffffff",
   55365 => x"ffffff",
   55366 => x"ffffff",
   55367 => x"ffffff",
   55368 => x"ffffff",
   55369 => x"ffffff",
   55370 => x"ffffff",
   55371 => x"ffffff",
   55372 => x"ffffff",
   55373 => x"ffffff",
   55374 => x"ffffff",
   55375 => x"ffffff",
   55376 => x"ffffff",
   55377 => x"ffffff",
   55378 => x"ffffff",
   55379 => x"ffffff",
   55380 => x"ffffff",
   55381 => x"ffffff",
   55382 => x"ffffff",
   55383 => x"ffffff",
   55384 => x"ffffff",
   55385 => x"ffffff",
   55386 => x"ffffff",
   55387 => x"ffffff",
   55388 => x"ffffff",
   55389 => x"ffffff",
   55390 => x"ffffff",
   55391 => x"ffffff",
   55392 => x"ffffff",
   55393 => x"ffffff",
   55394 => x"ffffff",
   55395 => x"ffffff",
   55396 => x"ffffff",
   55397 => x"ffffff",
   55398 => x"ffffff",
   55399 => x"ffffff",
   55400 => x"ffffff",
   55401 => x"ffffff",
   55402 => x"ffffff",
   55403 => x"ffffff",
   55404 => x"ffffff",
   55405 => x"ffffff",
   55406 => x"ffffff",
   55407 => x"ffffff",
   55408 => x"ffffff",
   55409 => x"ffffff",
   55410 => x"ffffff",
   55411 => x"ffffff",
   55412 => x"ffffff",
   55413 => x"ffffff",
   55414 => x"ffffff",
   55415 => x"ffffff",
   55416 => x"ffffff",
   55417 => x"ffffff",
   55418 => x"ffffff",
   55419 => x"ffffff",
   55420 => x"ffffff",
   55421 => x"ffffff",
   55422 => x"ffffff",
   55423 => x"ffffff",
   55424 => x"ffffff",
   55425 => x"ffffff",
   55426 => x"ffffff",
   55427 => x"ffffff",
   55428 => x"ffffff",
   55429 => x"fffa95",
   55430 => x"abffff",
   55431 => x"ffffff",
   55432 => x"ffffff",
   55433 => x"ffffff",
   55434 => x"ffffff",
   55435 => x"ffffff",
   55436 => x"ffffff",
   55437 => x"ffffff",
   55438 => x"ffffff",
   55439 => x"ffffff",
   55440 => x"ffffff",
   55441 => x"fffac3",
   55442 => x"0c30c3",
   55443 => x"0c30c3",
   55444 => x"0c30c3",
   55445 => x"0c30c3",
   55446 => x"0c30c3",
   55447 => x"0c30c3",
   55448 => x"0c30c3",
   55449 => x"0c30c3",
   55450 => x"0c30c3",
   55451 => x"0c30c3",
   55452 => x"0c30c3",
   55453 => x"082082",
   55454 => x"082082",
   55455 => x"082082",
   55456 => x"082082",
   55457 => x"082082",
   55458 => x"082082",
   55459 => x"082082",
   55460 => x"082082",
   55461 => x"082082",
   55462 => x"082082",
   55463 => x"082082",
   55464 => x"082082",
   55465 => x"082082",
   55466 => x"082082",
   55467 => x"082082",
   55468 => x"082082",
   55469 => x"082082",
   55470 => x"082082",
   55471 => x"082082",
   55472 => x"082082",
   55473 => x"082082",
   55474 => x"082082",
   55475 => x"082041",
   55476 => x"041041",
   55477 => x"041041",
   55478 => x"041041",
   55479 => x"041041",
   55480 => x"041041",
   55481 => x"041041",
   55482 => x"041041",
   55483 => x"041041",
   55484 => x"041041",
   55485 => x"041041",
   55486 => x"041041",
   55487 => x"041041",
   55488 => x"041041",
   55489 => x"041041",
   55490 => x"041041",
   55491 => x"041041",
   55492 => x"041041",
   55493 => x"041041",
   55494 => x"041041",
   55495 => x"041041",
   55496 => x"041041",
   55497 => x"041041",
   55498 => x"041000",
   55499 => x"000000",
   55500 => x"000000",
   55501 => x"000000",
   55502 => x"000000",
   55503 => x"000000",
   55504 => x"000000",
   55505 => x"000000",
   55506 => x"000000",
   55507 => x"000000",
   55508 => x"000000",
   55509 => x"00057f",
   55510 => x"ffffff",
   55511 => x"ffffff",
   55512 => x"ffffff",
   55513 => x"ffffd5",
   55514 => x"00002a",
   55515 => x"ffffff",
   55516 => x"ffffff",
   55517 => x"fff540",
   55518 => x"000015",
   55519 => x"ffffff",
   55520 => x"ffffff",
   55521 => x"ffffff",
   55522 => x"ffffff",
   55523 => x"ffffff",
   55524 => x"ffffff",
   55525 => x"ffffff",
   55526 => x"ffffff",
   55527 => x"ffffff",
   55528 => x"ffffff",
   55529 => x"ffffff",
   55530 => x"ffffff",
   55531 => x"ffffff",
   55532 => x"ffffff",
   55533 => x"ffffff",
   55534 => x"ffffff",
   55535 => x"ffffff",
   55536 => x"ffffff",
   55537 => x"ffffff",
   55538 => x"ffffff",
   55539 => x"ffffff",
   55540 => x"ffffff",
   55541 => x"ffffff",
   55542 => x"ffffff",
   55543 => x"ffffff",
   55544 => x"ffffff",
   55545 => x"ffffff",
   55546 => x"ffffff",
   55547 => x"ffffff",
   55548 => x"ffffff",
   55549 => x"ffffff",
   55550 => x"ffffff",
   55551 => x"ffffff",
   55552 => x"ffffff",
   55553 => x"ffffff",
   55554 => x"ffffff",
   55555 => x"ffffff",
   55556 => x"ffffff",
   55557 => x"ffffff",
   55558 => x"ffffff",
   55559 => x"ffffff",
   55560 => x"ffffff",
   55561 => x"ffffff",
   55562 => x"ffffff",
   55563 => x"ffffff",
   55564 => x"ffffff",
   55565 => x"ffffff",
   55566 => x"ffffff",
   55567 => x"ffffff",
   55568 => x"ffffff",
   55569 => x"ffffff",
   55570 => x"ffffff",
   55571 => x"ffffff",
   55572 => x"ffffff",
   55573 => x"ffffff",
   55574 => x"ffffff",
   55575 => x"ffffff",
   55576 => x"ffffff",
   55577 => x"ffffff",
   55578 => x"ffffff",
   55579 => x"ffffff",
   55580 => x"ffffff",
   55581 => x"ffffff",
   55582 => x"ffffff",
   55583 => x"ffffff",
   55584 => x"ffffff",
   55585 => x"ffffff",
   55586 => x"ffffff",
   55587 => x"ffffff",
   55588 => x"ffffff",
   55589 => x"fffa95",
   55590 => x"abffff",
   55591 => x"ffffff",
   55592 => x"ffffff",
   55593 => x"ffffff",
   55594 => x"ffffff",
   55595 => x"ffffff",
   55596 => x"ffffff",
   55597 => x"ffffff",
   55598 => x"ffffff",
   55599 => x"ffffff",
   55600 => x"ffffff",
   55601 => x"fffac3",
   55602 => x"0c30c3",
   55603 => x"0c30c3",
   55604 => x"0c30c3",
   55605 => x"0c30c3",
   55606 => x"0c30c3",
   55607 => x"0c30c3",
   55608 => x"0c30c3",
   55609 => x"0c30c3",
   55610 => x"0c30c3",
   55611 => x"0c30c3",
   55612 => x"0c30c3",
   55613 => x"082082",
   55614 => x"082082",
   55615 => x"082082",
   55616 => x"082082",
   55617 => x"082082",
   55618 => x"082082",
   55619 => x"082082",
   55620 => x"082082",
   55621 => x"082082",
   55622 => x"082082",
   55623 => x"082082",
   55624 => x"082082",
   55625 => x"082082",
   55626 => x"082082",
   55627 => x"082082",
   55628 => x"082082",
   55629 => x"082082",
   55630 => x"082082",
   55631 => x"082082",
   55632 => x"082082",
   55633 => x"082082",
   55634 => x"082082",
   55635 => x"082041",
   55636 => x"041041",
   55637 => x"041041",
   55638 => x"041041",
   55639 => x"041041",
   55640 => x"041041",
   55641 => x"041041",
   55642 => x"041041",
   55643 => x"041041",
   55644 => x"041041",
   55645 => x"041041",
   55646 => x"041041",
   55647 => x"041041",
   55648 => x"041041",
   55649 => x"041041",
   55650 => x"041041",
   55651 => x"041041",
   55652 => x"041041",
   55653 => x"041041",
   55654 => x"041041",
   55655 => x"041041",
   55656 => x"041041",
   55657 => x"041041",
   55658 => x"041000",
   55659 => x"000000",
   55660 => x"000000",
   55661 => x"000000",
   55662 => x"000000",
   55663 => x"000000",
   55664 => x"000000",
   55665 => x"000000",
   55666 => x"000000",
   55667 => x"000000",
   55668 => x"000000",
   55669 => x"00057f",
   55670 => x"ffffff",
   55671 => x"ffffff",
   55672 => x"ffffff",
   55673 => x"ffffd5",
   55674 => x"000015",
   55675 => x"aaaaaa",
   55676 => x"aaaa95",
   55677 => x"555000",
   55678 => x"00002a",
   55679 => x"ffffff",
   55680 => x"ffffff",
   55681 => x"ffffff",
   55682 => x"ffffff",
   55683 => x"ffffff",
   55684 => x"ffffff",
   55685 => x"ffffff",
   55686 => x"ffffff",
   55687 => x"ffffff",
   55688 => x"ffffff",
   55689 => x"ffffff",
   55690 => x"ffffff",
   55691 => x"ffffff",
   55692 => x"ffffff",
   55693 => x"ffffff",
   55694 => x"ffffff",
   55695 => x"ffffff",
   55696 => x"ffffff",
   55697 => x"ffffff",
   55698 => x"ffffff",
   55699 => x"ffffff",
   55700 => x"ffffff",
   55701 => x"ffffff",
   55702 => x"ffffff",
   55703 => x"ffffff",
   55704 => x"ffffff",
   55705 => x"ffffff",
   55706 => x"ffffff",
   55707 => x"ffffff",
   55708 => x"ffffff",
   55709 => x"ffffff",
   55710 => x"ffffff",
   55711 => x"ffffff",
   55712 => x"ffffff",
   55713 => x"ffffff",
   55714 => x"ffffff",
   55715 => x"ffffff",
   55716 => x"ffffff",
   55717 => x"ffffff",
   55718 => x"ffffff",
   55719 => x"ffffff",
   55720 => x"ffffff",
   55721 => x"ffffff",
   55722 => x"ffffff",
   55723 => x"ffffff",
   55724 => x"ffffff",
   55725 => x"ffffff",
   55726 => x"ffffff",
   55727 => x"ffffff",
   55728 => x"ffffff",
   55729 => x"ffffff",
   55730 => x"ffffff",
   55731 => x"ffffff",
   55732 => x"ffffff",
   55733 => x"ffffff",
   55734 => x"ffffff",
   55735 => x"ffffff",
   55736 => x"ffffff",
   55737 => x"ffffff",
   55738 => x"ffffff",
   55739 => x"ffffff",
   55740 => x"ffffff",
   55741 => x"ffffff",
   55742 => x"ffffff",
   55743 => x"ffffff",
   55744 => x"ffffff",
   55745 => x"ffffff",
   55746 => x"ffffff",
   55747 => x"ffffff",
   55748 => x"ffffff",
   55749 => x"fffa95",
   55750 => x"abffff",
   55751 => x"ffffff",
   55752 => x"ffffff",
   55753 => x"ffffff",
   55754 => x"ffffff",
   55755 => x"ffffff",
   55756 => x"ffffff",
   55757 => x"ffffff",
   55758 => x"ffffff",
   55759 => x"ffffff",
   55760 => x"ffffff",
   55761 => x"fffac3",
   55762 => x"0c30c3",
   55763 => x"0c30c3",
   55764 => x"0c30c3",
   55765 => x"0c30c3",
   55766 => x"0c30c3",
   55767 => x"0c30c3",
   55768 => x"0c30c3",
   55769 => x"0c30c3",
   55770 => x"0c30c3",
   55771 => x"0c30c3",
   55772 => x"0c30c3",
   55773 => x"082082",
   55774 => x"082082",
   55775 => x"082082",
   55776 => x"082082",
   55777 => x"082082",
   55778 => x"082082",
   55779 => x"082082",
   55780 => x"082082",
   55781 => x"082082",
   55782 => x"082082",
   55783 => x"082082",
   55784 => x"082082",
   55785 => x"082082",
   55786 => x"082082",
   55787 => x"082082",
   55788 => x"082082",
   55789 => x"082082",
   55790 => x"082082",
   55791 => x"082082",
   55792 => x"082082",
   55793 => x"082082",
   55794 => x"082082",
   55795 => x"082041",
   55796 => x"041041",
   55797 => x"041041",
   55798 => x"041041",
   55799 => x"041041",
   55800 => x"041041",
   55801 => x"041041",
   55802 => x"041041",
   55803 => x"041041",
   55804 => x"041041",
   55805 => x"041041",
   55806 => x"041041",
   55807 => x"041041",
   55808 => x"041041",
   55809 => x"041041",
   55810 => x"041041",
   55811 => x"041041",
   55812 => x"041041",
   55813 => x"041041",
   55814 => x"041041",
   55815 => x"041041",
   55816 => x"041041",
   55817 => x"041041",
   55818 => x"041000",
   55819 => x"000000",
   55820 => x"000000",
   55821 => x"000000",
   55822 => x"000000",
   55823 => x"000000",
   55824 => x"000000",
   55825 => x"000000",
   55826 => x"000000",
   55827 => x"000000",
   55828 => x"000000",
   55829 => x"00057f",
   55830 => x"ffffff",
   55831 => x"ffffff",
   55832 => x"ffffff",
   55833 => x"ffffd5",
   55834 => x"000000",
   55835 => x"000000",
   55836 => x"000000",
   55837 => x"000000",
   55838 => x"000abf",
   55839 => x"ffffff",
   55840 => x"ffffff",
   55841 => x"ffffff",
   55842 => x"ffffff",
   55843 => x"ffffff",
   55844 => x"ffffff",
   55845 => x"ffffff",
   55846 => x"ffffff",
   55847 => x"ffffff",
   55848 => x"ffffff",
   55849 => x"ffffff",
   55850 => x"ffffff",
   55851 => x"ffffff",
   55852 => x"ffffff",
   55853 => x"ffffff",
   55854 => x"ffffff",
   55855 => x"ffffff",
   55856 => x"ffffff",
   55857 => x"ffffff",
   55858 => x"ffffff",
   55859 => x"ffffff",
   55860 => x"ffffff",
   55861 => x"ffffff",
   55862 => x"ffffff",
   55863 => x"ffffff",
   55864 => x"ffffff",
   55865 => x"ffffff",
   55866 => x"ffffff",
   55867 => x"ffffff",
   55868 => x"ffffff",
   55869 => x"ffffff",
   55870 => x"ffffff",
   55871 => x"ffffff",
   55872 => x"ffffff",
   55873 => x"ffffff",
   55874 => x"ffffff",
   55875 => x"ffffff",
   55876 => x"ffffff",
   55877 => x"ffffff",
   55878 => x"ffffff",
   55879 => x"ffffff",
   55880 => x"ffffff",
   55881 => x"ffffff",
   55882 => x"ffffff",
   55883 => x"ffffff",
   55884 => x"ffffff",
   55885 => x"ffffff",
   55886 => x"ffffff",
   55887 => x"ffffff",
   55888 => x"ffffff",
   55889 => x"ffffff",
   55890 => x"ffffff",
   55891 => x"ffffff",
   55892 => x"ffffff",
   55893 => x"ffffff",
   55894 => x"ffffff",
   55895 => x"ffffff",
   55896 => x"ffffff",
   55897 => x"ffffff",
   55898 => x"ffffff",
   55899 => x"ffffff",
   55900 => x"ffffff",
   55901 => x"ffffff",
   55902 => x"ffffff",
   55903 => x"ffffff",
   55904 => x"ffffff",
   55905 => x"ffffff",
   55906 => x"ffffff",
   55907 => x"ffffff",
   55908 => x"ffffff",
   55909 => x"fffa95",
   55910 => x"abffff",
   55911 => x"ffffff",
   55912 => x"ffffff",
   55913 => x"ffffff",
   55914 => x"ffffff",
   55915 => x"ffffff",
   55916 => x"ffffff",
   55917 => x"ffffff",
   55918 => x"ffffff",
   55919 => x"ffffff",
   55920 => x"ffffff",
   55921 => x"fffac3",
   55922 => x"0c30c3",
   55923 => x"0c30c3",
   55924 => x"0c30c3",
   55925 => x"0c30c3",
   55926 => x"0c30c3",
   55927 => x"0c30c3",
   55928 => x"0c30c3",
   55929 => x"0c30c3",
   55930 => x"0c30c3",
   55931 => x"0c30c3",
   55932 => x"0c30c3",
   55933 => x"082082",
   55934 => x"082082",
   55935 => x"082082",
   55936 => x"082082",
   55937 => x"082082",
   55938 => x"082082",
   55939 => x"082082",
   55940 => x"082082",
   55941 => x"082082",
   55942 => x"082082",
   55943 => x"082082",
   55944 => x"082082",
   55945 => x"082082",
   55946 => x"082082",
   55947 => x"082082",
   55948 => x"082082",
   55949 => x"082082",
   55950 => x"082082",
   55951 => x"082082",
   55952 => x"082082",
   55953 => x"082082",
   55954 => x"082082",
   55955 => x"082041",
   55956 => x"041041",
   55957 => x"041041",
   55958 => x"041041",
   55959 => x"041041",
   55960 => x"041041",
   55961 => x"041041",
   55962 => x"041041",
   55963 => x"041041",
   55964 => x"041041",
   55965 => x"041041",
   55966 => x"041041",
   55967 => x"041041",
   55968 => x"041041",
   55969 => x"041041",
   55970 => x"041041",
   55971 => x"041041",
   55972 => x"041041",
   55973 => x"041041",
   55974 => x"041041",
   55975 => x"041041",
   55976 => x"041041",
   55977 => x"041041",
   55978 => x"041000",
   55979 => x"000000",
   55980 => x"000000",
   55981 => x"000000",
   55982 => x"000000",
   55983 => x"000000",
   55984 => x"000000",
   55985 => x"000000",
   55986 => x"000000",
   55987 => x"000000",
   55988 => x"000000",
   55989 => x"00057f",
   55990 => x"ffffff",
   55991 => x"ffffff",
   55992 => x"ffffff",
   55993 => x"ffffd5",
   55994 => x"000000",
   55995 => x"000000",
   55996 => x"000000",
   55997 => x"000000",
   55998 => x"56afff",
   55999 => x"ffffff",
   56000 => x"ffffff",
   56001 => x"ffffff",
   56002 => x"ffffff",
   56003 => x"ffffff",
   56004 => x"ffffff",
   56005 => x"ffffff",
   56006 => x"ffffff",
   56007 => x"ffffff",
   56008 => x"ffffff",
   56009 => x"ffffff",
   56010 => x"ffffff",
   56011 => x"ffffff",
   56012 => x"ffffff",
   56013 => x"ffffff",
   56014 => x"ffffff",
   56015 => x"ffffff",
   56016 => x"ffffff",
   56017 => x"ffffff",
   56018 => x"ffffff",
   56019 => x"ffffff",
   56020 => x"ffffff",
   56021 => x"ffffff",
   56022 => x"ffffff",
   56023 => x"ffffff",
   56024 => x"ffffff",
   56025 => x"ffffff",
   56026 => x"ffffff",
   56027 => x"ffffff",
   56028 => x"ffffff",
   56029 => x"ffffff",
   56030 => x"ffffff",
   56031 => x"ffffff",
   56032 => x"ffffff",
   56033 => x"ffffff",
   56034 => x"ffffff",
   56035 => x"ffffff",
   56036 => x"ffffff",
   56037 => x"ffffff",
   56038 => x"ffffff",
   56039 => x"ffffff",
   56040 => x"ffffff",
   56041 => x"ffffff",
   56042 => x"ffffff",
   56043 => x"ffffff",
   56044 => x"ffffff",
   56045 => x"ffffff",
   56046 => x"ffffff",
   56047 => x"ffffff",
   56048 => x"ffffff",
   56049 => x"ffffff",
   56050 => x"ffffff",
   56051 => x"ffffff",
   56052 => x"ffffff",
   56053 => x"ffffff",
   56054 => x"ffffff",
   56055 => x"ffffff",
   56056 => x"ffffff",
   56057 => x"ffffff",
   56058 => x"ffffff",
   56059 => x"ffffff",
   56060 => x"ffffff",
   56061 => x"ffffff",
   56062 => x"ffffff",
   56063 => x"ffffff",
   56064 => x"ffffff",
   56065 => x"ffffff",
   56066 => x"ffffff",
   56067 => x"ffffff",
   56068 => x"ffffff",
   56069 => x"fffa95",
   56070 => x"abffff",
   56071 => x"ffffff",
   56072 => x"ffffff",
   56073 => x"ffffff",
   56074 => x"ffffff",
   56075 => x"ffffff",
   56076 => x"ffffff",
   56077 => x"ffffff",
   56078 => x"ffffff",
   56079 => x"ffffff",
   56080 => x"ffffff",
   56081 => x"fffac3",
   56082 => x"0c30c3",
   56083 => x"0c30c3",
   56084 => x"0c30c3",
   56085 => x"0c30c3",
   56086 => x"0c30c3",
   56087 => x"0c30c3",
   56088 => x"0c30c3",
   56089 => x"0c30c3",
   56090 => x"0c30c3",
   56091 => x"0c30c3",
   56092 => x"0c30c3",
   56093 => x"082082",
   56094 => x"082082",
   56095 => x"082082",
   56096 => x"082082",
   56097 => x"082082",
   56098 => x"082082",
   56099 => x"082082",
   56100 => x"082082",
   56101 => x"082082",
   56102 => x"082082",
   56103 => x"082082",
   56104 => x"082082",
   56105 => x"082082",
   56106 => x"082082",
   56107 => x"082082",
   56108 => x"082082",
   56109 => x"082082",
   56110 => x"082082",
   56111 => x"082082",
   56112 => x"082082",
   56113 => x"082082",
   56114 => x"082082",
   56115 => x"082041",
   56116 => x"041041",
   56117 => x"041041",
   56118 => x"041041",
   56119 => x"041041",
   56120 => x"041041",
   56121 => x"041041",
   56122 => x"041041",
   56123 => x"041041",
   56124 => x"041041",
   56125 => x"041041",
   56126 => x"041041",
   56127 => x"041041",
   56128 => x"041041",
   56129 => x"041041",
   56130 => x"041041",
   56131 => x"041041",
   56132 => x"041041",
   56133 => x"041041",
   56134 => x"041041",
   56135 => x"041041",
   56136 => x"041041",
   56137 => x"041041",
   56138 => x"041000",
   56139 => x"000000",
   56140 => x"000000",
   56141 => x"000000",
   56142 => x"000000",
   56143 => x"000000",
   56144 => x"000000",
   56145 => x"000000",
   56146 => x"000000",
   56147 => x"000000",
   56148 => x"000000",
   56149 => x"00057f",
   56150 => x"ffffff",
   56151 => x"ffffff",
   56152 => x"ffffff",
   56153 => x"ffffd5",
   56154 => x"000000",
   56155 => x"000000",
   56156 => x"000015",
   56157 => x"555aaa",
   56158 => x"ffffff",
   56159 => x"ffffff",
   56160 => x"ffffff",
   56161 => x"ffffff",
   56162 => x"ffffff",
   56163 => x"ffffff",
   56164 => x"ffffff",
   56165 => x"ffffff",
   56166 => x"ffffff",
   56167 => x"ffffff",
   56168 => x"ffffff",
   56169 => x"ffffff",
   56170 => x"ffffff",
   56171 => x"ffffff",
   56172 => x"ffffff",
   56173 => x"ffffff",
   56174 => x"ffffff",
   56175 => x"ffffff",
   56176 => x"ffffff",
   56177 => x"ffffff",
   56178 => x"ffffff",
   56179 => x"ffffff",
   56180 => x"ffffff",
   56181 => x"ffffff",
   56182 => x"ffffff",
   56183 => x"ffffff",
   56184 => x"ffffff",
   56185 => x"ffffff",
   56186 => x"ffffff",
   56187 => x"ffffff",
   56188 => x"ffffff",
   56189 => x"ffffff",
   56190 => x"ffffff",
   56191 => x"ffffff",
   56192 => x"ffffff",
   56193 => x"ffffff",
   56194 => x"ffffff",
   56195 => x"ffffff",
   56196 => x"ffffff",
   56197 => x"ffffff",
   56198 => x"ffffff",
   56199 => x"ffffff",
   56200 => x"ffffff",
   56201 => x"ffffff",
   56202 => x"ffffff",
   56203 => x"ffffff",
   56204 => x"ffffff",
   56205 => x"ffffff",
   56206 => x"ffffff",
   56207 => x"ffffff",
   56208 => x"ffffff",
   56209 => x"ffffff",
   56210 => x"ffffff",
   56211 => x"ffffff",
   56212 => x"ffffff",
   56213 => x"ffffff",
   56214 => x"ffffff",
   56215 => x"ffffff",
   56216 => x"ffffff",
   56217 => x"ffffff",
   56218 => x"ffffff",
   56219 => x"ffffff",
   56220 => x"ffffff",
   56221 => x"ffffff",
   56222 => x"ffffff",
   56223 => x"ffffff",
   56224 => x"ffffff",
   56225 => x"ffffff",
   56226 => x"ffffff",
   56227 => x"ffffff",
   56228 => x"ffffff",
   56229 => x"fffa95",
   56230 => x"abffff",
   56231 => x"ffffff",
   56232 => x"ffffff",
   56233 => x"ffffff",
   56234 => x"ffffff",
   56235 => x"ffffff",
   56236 => x"ffffff",
   56237 => x"ffffff",
   56238 => x"ffffff",
   56239 => x"ffffff",
   56240 => x"ffffff",
   56241 => x"fffac3",
   56242 => x"0c30c3",
   56243 => x"0c30c3",
   56244 => x"0c30c3",
   56245 => x"0c30c3",
   56246 => x"0c30c3",
   56247 => x"0c30c3",
   56248 => x"0c30c3",
   56249 => x"0c30c3",
   56250 => x"0c30c3",
   56251 => x"0c30c3",
   56252 => x"0c30c3",
   56253 => x"082082",
   56254 => x"082082",
   56255 => x"082082",
   56256 => x"082082",
   56257 => x"082082",
   56258 => x"082082",
   56259 => x"082082",
   56260 => x"082082",
   56261 => x"082082",
   56262 => x"082082",
   56263 => x"082082",
   56264 => x"082082",
   56265 => x"082082",
   56266 => x"082082",
   56267 => x"082082",
   56268 => x"082082",
   56269 => x"082082",
   56270 => x"082082",
   56271 => x"082082",
   56272 => x"082082",
   56273 => x"082082",
   56274 => x"082082",
   56275 => x"082041",
   56276 => x"041041",
   56277 => x"041041",
   56278 => x"041041",
   56279 => x"041041",
   56280 => x"041041",
   56281 => x"041041",
   56282 => x"041041",
   56283 => x"041041",
   56284 => x"041041",
   56285 => x"041041",
   56286 => x"041041",
   56287 => x"041041",
   56288 => x"041041",
   56289 => x"041041",
   56290 => x"041041",
   56291 => x"041041",
   56292 => x"041041",
   56293 => x"041041",
   56294 => x"041041",
   56295 => x"041041",
   56296 => x"041041",
   56297 => x"041041",
   56298 => x"041000",
   56299 => x"000000",
   56300 => x"000000",
   56301 => x"000000",
   56302 => x"000000",
   56303 => x"000000",
   56304 => x"000000",
   56305 => x"000000",
   56306 => x"000000",
   56307 => x"000000",
   56308 => x"000000",
   56309 => x"00057f",
   56310 => x"ffffff",
   56311 => x"ffffff",
   56312 => x"ffffff",
   56313 => x"ffffea",
   56314 => x"aaaaaa",
   56315 => x"aaaaaa",
   56316 => x"aaaaaa",
   56317 => x"abffff",
   56318 => x"ffffff",
   56319 => x"ffffff",
   56320 => x"ffffff",
   56321 => x"ffffff",
   56322 => x"ffffff",
   56323 => x"ffffff",
   56324 => x"ffffff",
   56325 => x"ffffff",
   56326 => x"ffffff",
   56327 => x"ffffff",
   56328 => x"ffffff",
   56329 => x"ffffff",
   56330 => x"ffffff",
   56331 => x"ffffff",
   56332 => x"ffffff",
   56333 => x"ffffff",
   56334 => x"ffffff",
   56335 => x"ffffff",
   56336 => x"ffffff",
   56337 => x"ffffff",
   56338 => x"ffffff",
   56339 => x"ffffff",
   56340 => x"ffffff",
   56341 => x"ffffff",
   56342 => x"ffffff",
   56343 => x"ffffff",
   56344 => x"ffffff",
   56345 => x"ffffff",
   56346 => x"ffffff",
   56347 => x"ffffff",
   56348 => x"ffffff",
   56349 => x"ffffff",
   56350 => x"ffffff",
   56351 => x"ffffff",
   56352 => x"ffffff",
   56353 => x"ffffff",
   56354 => x"ffffff",
   56355 => x"ffffff",
   56356 => x"ffffff",
   56357 => x"ffffff",
   56358 => x"ffffff",
   56359 => x"ffffff",
   56360 => x"ffffff",
   56361 => x"ffffff",
   56362 => x"ffffff",
   56363 => x"ffffff",
   56364 => x"ffffff",
   56365 => x"ffffff",
   56366 => x"ffffff",
   56367 => x"ffffff",
   56368 => x"ffffff",
   56369 => x"ffffff",
   56370 => x"ffffff",
   56371 => x"ffffff",
   56372 => x"ffffff",
   56373 => x"ffffff",
   56374 => x"ffffff",
   56375 => x"ffffff",
   56376 => x"ffffff",
   56377 => x"ffffff",
   56378 => x"ffffff",
   56379 => x"ffffff",
   56380 => x"ffffff",
   56381 => x"ffffff",
   56382 => x"ffffff",
   56383 => x"ffffff",
   56384 => x"ffffff",
   56385 => x"ffffff",
   56386 => x"ffffff",
   56387 => x"ffffff",
   56388 => x"ffffff",
   56389 => x"fffa95",
   56390 => x"abffff",
   56391 => x"ffffff",
   56392 => x"ffffff",
   56393 => x"ffffff",
   56394 => x"ffffff",
   56395 => x"ffffff",
   56396 => x"ffffff",
   56397 => x"ffffff",
   56398 => x"ffffff",
   56399 => x"ffffff",
   56400 => x"ffffff",
   56401 => x"fffac3",
   56402 => x"0c30c3",
   56403 => x"0c30c3",
   56404 => x"0c30c3",
   56405 => x"0c30c3",
   56406 => x"0c30c3",
   56407 => x"0c30c3",
   56408 => x"0c30c3",
   56409 => x"0c30c3",
   56410 => x"0c30c3",
   56411 => x"0c30c3",
   56412 => x"0c30c3",
   56413 => x"082082",
   56414 => x"082082",
   56415 => x"082082",
   56416 => x"082082",
   56417 => x"082082",
   56418 => x"082082",
   56419 => x"082082",
   56420 => x"082082",
   56421 => x"082082",
   56422 => x"082082",
   56423 => x"082082",
   56424 => x"082082",
   56425 => x"082082",
   56426 => x"082082",
   56427 => x"082082",
   56428 => x"082082",
   56429 => x"082082",
   56430 => x"082082",
   56431 => x"082082",
   56432 => x"082082",
   56433 => x"082082",
   56434 => x"082082",
   56435 => x"082041",
   56436 => x"041041",
   56437 => x"041041",
   56438 => x"041041",
   56439 => x"041041",
   56440 => x"041041",
   56441 => x"041041",
   56442 => x"041041",
   56443 => x"041041",
   56444 => x"041041",
   56445 => x"041041",
   56446 => x"041041",
   56447 => x"041041",
   56448 => x"041041",
   56449 => x"041041",
   56450 => x"041041",
   56451 => x"041041",
   56452 => x"041041",
   56453 => x"041041",
   56454 => x"041041",
   56455 => x"041041",
   56456 => x"041041",
   56457 => x"041041",
   56458 => x"041000",
   56459 => x"000000",
   56460 => x"000000",
   56461 => x"000000",
   56462 => x"000000",
   56463 => x"000000",
   56464 => x"000000",
   56465 => x"000000",
   56466 => x"000000",
   56467 => x"000000",
   56468 => x"000000",
   56469 => x"00057f",
   56470 => x"ffffff",
   56471 => x"ffffff",
   56472 => x"ffffff",
   56473 => x"ffffff",
   56474 => x"ffffff",
   56475 => x"ffffff",
   56476 => x"ffffff",
   56477 => x"ffffff",
   56478 => x"ffffff",
   56479 => x"ffffff",
   56480 => x"ffffff",
   56481 => x"ffffff",
   56482 => x"ffffff",
   56483 => x"ffffff",
   56484 => x"ffffff",
   56485 => x"ffffff",
   56486 => x"ffffff",
   56487 => x"ffffff",
   56488 => x"ffffff",
   56489 => x"ffffff",
   56490 => x"ffffff",
   56491 => x"ffffff",
   56492 => x"ffffff",
   56493 => x"ffffff",
   56494 => x"ffffff",
   56495 => x"ffffff",
   56496 => x"ffffff",
   56497 => x"ffffff",
   56498 => x"ffffff",
   56499 => x"ffffff",
   56500 => x"ffffff",
   56501 => x"ffffff",
   56502 => x"ffffff",
   56503 => x"ffffff",
   56504 => x"ffffff",
   56505 => x"ffffff",
   56506 => x"ffffff",
   56507 => x"ffffff",
   56508 => x"ffffff",
   56509 => x"ffffff",
   56510 => x"ffffff",
   56511 => x"ffffff",
   56512 => x"ffffff",
   56513 => x"ffffff",
   56514 => x"ffffff",
   56515 => x"ffffff",
   56516 => x"ffffff",
   56517 => x"ffffff",
   56518 => x"ffffff",
   56519 => x"ffffff",
   56520 => x"ffffff",
   56521 => x"ffffff",
   56522 => x"ffffff",
   56523 => x"ffffff",
   56524 => x"ffffff",
   56525 => x"ffffff",
   56526 => x"ffffff",
   56527 => x"ffffff",
   56528 => x"ffffff",
   56529 => x"ffffff",
   56530 => x"ffffff",
   56531 => x"ffffff",
   56532 => x"ffffff",
   56533 => x"ffffff",
   56534 => x"ffffff",
   56535 => x"ffffff",
   56536 => x"ffffff",
   56537 => x"ffffff",
   56538 => x"ffffff",
   56539 => x"ffffff",
   56540 => x"ffffff",
   56541 => x"ffffff",
   56542 => x"ffffff",
   56543 => x"ffffff",
   56544 => x"ffffff",
   56545 => x"ffffff",
   56546 => x"ffffff",
   56547 => x"ffffff",
   56548 => x"ffffff",
   56549 => x"fffa95",
   56550 => x"abffff",
   56551 => x"ffffff",
   56552 => x"ffffff",
   56553 => x"ffffff",
   56554 => x"ffffff",
   56555 => x"ffffff",
   56556 => x"ffffff",
   56557 => x"ffffff",
   56558 => x"ffffff",
   56559 => x"ffffff",
   56560 => x"ffffff",
   56561 => x"fffac3",
   56562 => x"0c30c3",
   56563 => x"0c30c3",
   56564 => x"0c30c3",
   56565 => x"0c30c3",
   56566 => x"0c30c3",
   56567 => x"0c30c3",
   56568 => x"0c30c3",
   56569 => x"0c30c3",
   56570 => x"0c30c3",
   56571 => x"0c30c3",
   56572 => x"0c30c3",
   56573 => x"082082",
   56574 => x"082082",
   56575 => x"082082",
   56576 => x"082082",
   56577 => x"082082",
   56578 => x"082082",
   56579 => x"082082",
   56580 => x"082082",
   56581 => x"082082",
   56582 => x"082082",
   56583 => x"082082",
   56584 => x"082082",
   56585 => x"082082",
   56586 => x"082082",
   56587 => x"082082",
   56588 => x"082082",
   56589 => x"082082",
   56590 => x"082082",
   56591 => x"082082",
   56592 => x"082082",
   56593 => x"082082",
   56594 => x"082082",
   56595 => x"082041",
   56596 => x"041041",
   56597 => x"041041",
   56598 => x"041041",
   56599 => x"041041",
   56600 => x"041041",
   56601 => x"041041",
   56602 => x"041041",
   56603 => x"041041",
   56604 => x"041041",
   56605 => x"041041",
   56606 => x"041041",
   56607 => x"041041",
   56608 => x"041041",
   56609 => x"041041",
   56610 => x"041041",
   56611 => x"041041",
   56612 => x"041041",
   56613 => x"041041",
   56614 => x"041041",
   56615 => x"041041",
   56616 => x"041041",
   56617 => x"041041",
   56618 => x"041000",
   56619 => x"000000",
   56620 => x"000000",
   56621 => x"000000",
   56622 => x"000000",
   56623 => x"000000",
   56624 => x"000000",
   56625 => x"000000",
   56626 => x"000000",
   56627 => x"000000",
   56628 => x"000000",
   56629 => x"00057f",
   56630 => x"ffffff",
   56631 => x"ffffff",
   56632 => x"ffffff",
   56633 => x"ffffff",
   56634 => x"ffffff",
   56635 => x"ffffff",
   56636 => x"ffffff",
   56637 => x"ffffff",
   56638 => x"ffffff",
   56639 => x"ffffff",
   56640 => x"ffffff",
   56641 => x"ffffff",
   56642 => x"ffffff",
   56643 => x"ffffff",
   56644 => x"ffffff",
   56645 => x"ffffff",
   56646 => x"ffffff",
   56647 => x"ffffff",
   56648 => x"ffffff",
   56649 => x"ffffff",
   56650 => x"ffffff",
   56651 => x"ffffff",
   56652 => x"ffffff",
   56653 => x"ffffff",
   56654 => x"ffffff",
   56655 => x"ffffff",
   56656 => x"ffffff",
   56657 => x"ffffff",
   56658 => x"ffffff",
   56659 => x"ffffff",
   56660 => x"ffffff",
   56661 => x"ffffff",
   56662 => x"ffffff",
   56663 => x"ffffff",
   56664 => x"ffffff",
   56665 => x"ffffff",
   56666 => x"ffffff",
   56667 => x"ffffff",
   56668 => x"ffffff",
   56669 => x"ffffff",
   56670 => x"ffffff",
   56671 => x"ffffff",
   56672 => x"ffffff",
   56673 => x"ffffff",
   56674 => x"ffffff",
   56675 => x"ffffff",
   56676 => x"ffffff",
   56677 => x"ffffff",
   56678 => x"ffffff",
   56679 => x"ffffff",
   56680 => x"ffffff",
   56681 => x"ffffff",
   56682 => x"ffffff",
   56683 => x"ffffff",
   56684 => x"ffffff",
   56685 => x"ffffff",
   56686 => x"ffffff",
   56687 => x"ffffff",
   56688 => x"ffffff",
   56689 => x"ffffff",
   56690 => x"ffffff",
   56691 => x"ffffff",
   56692 => x"ffffff",
   56693 => x"ffffff",
   56694 => x"ffffff",
   56695 => x"ffffff",
   56696 => x"ffffff",
   56697 => x"ffffff",
   56698 => x"ffffff",
   56699 => x"ffffff",
   56700 => x"ffffff",
   56701 => x"ffffff",
   56702 => x"ffffff",
   56703 => x"ffffff",
   56704 => x"ffffff",
   56705 => x"ffffff",
   56706 => x"ffffff",
   56707 => x"ffffff",
   56708 => x"ffffff",
   56709 => x"fffa95",
   56710 => x"abffff",
   56711 => x"ffffff",
   56712 => x"ffffff",
   56713 => x"ffffff",
   56714 => x"ffffff",
   56715 => x"ffffff",
   56716 => x"ffffff",
   56717 => x"ffffff",
   56718 => x"ffffff",
   56719 => x"ffffff",
   56720 => x"ffffff",
   56721 => x"fffac3",
   56722 => x"0c30c3",
   56723 => x"0c30c3",
   56724 => x"0c30c3",
   56725 => x"0c30c3",
   56726 => x"0c30c3",
   56727 => x"0c30c3",
   56728 => x"0c30c3",
   56729 => x"0c30c3",
   56730 => x"0c30c3",
   56731 => x"0c30c3",
   56732 => x"0c30c3",
   56733 => x"082082",
   56734 => x"082082",
   56735 => x"082082",
   56736 => x"082082",
   56737 => x"082082",
   56738 => x"082082",
   56739 => x"082082",
   56740 => x"082082",
   56741 => x"082082",
   56742 => x"082082",
   56743 => x"082082",
   56744 => x"082082",
   56745 => x"082082",
   56746 => x"082082",
   56747 => x"082082",
   56748 => x"082082",
   56749 => x"082082",
   56750 => x"082082",
   56751 => x"082082",
   56752 => x"082082",
   56753 => x"082082",
   56754 => x"082082",
   56755 => x"082041",
   56756 => x"041041",
   56757 => x"041041",
   56758 => x"041041",
   56759 => x"041041",
   56760 => x"041041",
   56761 => x"041041",
   56762 => x"041041",
   56763 => x"041041",
   56764 => x"041041",
   56765 => x"041041",
   56766 => x"041041",
   56767 => x"041041",
   56768 => x"041041",
   56769 => x"041041",
   56770 => x"041041",
   56771 => x"041041",
   56772 => x"041041",
   56773 => x"041041",
   56774 => x"041041",
   56775 => x"041041",
   56776 => x"041041",
   56777 => x"041041",
   56778 => x"041000",
   56779 => x"000000",
   56780 => x"000000",
   56781 => x"000000",
   56782 => x"000000",
   56783 => x"000000",
   56784 => x"000000",
   56785 => x"000000",
   56786 => x"000000",
   56787 => x"000000",
   56788 => x"000000",
   56789 => x"00057f",
   56790 => x"ffffff",
   56791 => x"ffffff",
   56792 => x"ffffff",
   56793 => x"ffffff",
   56794 => x"ffffff",
   56795 => x"ffffff",
   56796 => x"ffffff",
   56797 => x"ffffff",
   56798 => x"ffffff",
   56799 => x"ffffff",
   56800 => x"ffffff",
   56801 => x"ffffff",
   56802 => x"ffffff",
   56803 => x"ffffff",
   56804 => x"ffffff",
   56805 => x"ffffff",
   56806 => x"ffffff",
   56807 => x"ffffff",
   56808 => x"ffffff",
   56809 => x"ffffff",
   56810 => x"ffffff",
   56811 => x"ffffff",
   56812 => x"ffffff",
   56813 => x"ffffff",
   56814 => x"ffffff",
   56815 => x"ffffff",
   56816 => x"ffffff",
   56817 => x"ffffff",
   56818 => x"ffffff",
   56819 => x"ffffff",
   56820 => x"ffffff",
   56821 => x"ffffff",
   56822 => x"ffffff",
   56823 => x"ffffff",
   56824 => x"ffffff",
   56825 => x"ffffff",
   56826 => x"ffffff",
   56827 => x"ffffff",
   56828 => x"ffffff",
   56829 => x"ffffff",
   56830 => x"ffffff",
   56831 => x"ffffff",
   56832 => x"ffffff",
   56833 => x"ffffff",
   56834 => x"ffffff",
   56835 => x"ffffff",
   56836 => x"ffffff",
   56837 => x"ffffff",
   56838 => x"ffffff",
   56839 => x"ffffff",
   56840 => x"ffffff",
   56841 => x"ffffff",
   56842 => x"ffffff",
   56843 => x"ffffff",
   56844 => x"ffffff",
   56845 => x"ffffff",
   56846 => x"ffffff",
   56847 => x"ffffff",
   56848 => x"ffffff",
   56849 => x"ffffff",
   56850 => x"ffffff",
   56851 => x"ffffff",
   56852 => x"ffffff",
   56853 => x"ffffff",
   56854 => x"ffffff",
   56855 => x"ffffff",
   56856 => x"ffffff",
   56857 => x"ffffff",
   56858 => x"ffffff",
   56859 => x"ffffff",
   56860 => x"ffffff",
   56861 => x"ffffff",
   56862 => x"ffffff",
   56863 => x"ffffff",
   56864 => x"ffffff",
   56865 => x"ffffff",
   56866 => x"ffffff",
   56867 => x"ffffff",
   56868 => x"ffffff",
   56869 => x"fffa95",
   56870 => x"abffff",
   56871 => x"ffffff",
   56872 => x"ffffff",
   56873 => x"ffffff",
   56874 => x"ffffff",
   56875 => x"ffffff",
   56876 => x"ffffff",
   56877 => x"ffffff",
   56878 => x"ffffff",
   56879 => x"ffffff",
   56880 => x"ffffff",
   56881 => x"fffac3",
   56882 => x"0c30c3",
   56883 => x"0c30c3",
   56884 => x"0c30c3",
   56885 => x"0c30c3",
   56886 => x"0c30c3",
   56887 => x"0c30c3",
   56888 => x"0c30c3",
   56889 => x"0c30c3",
   56890 => x"0c30c3",
   56891 => x"0c30c3",
   56892 => x"0c30c3",
   56893 => x"082082",
   56894 => x"082082",
   56895 => x"082082",
   56896 => x"082082",
   56897 => x"082082",
   56898 => x"082082",
   56899 => x"082082",
   56900 => x"082082",
   56901 => x"082082",
   56902 => x"082082",
   56903 => x"082082",
   56904 => x"082082",
   56905 => x"082082",
   56906 => x"082082",
   56907 => x"082082",
   56908 => x"082082",
   56909 => x"082082",
   56910 => x"082082",
   56911 => x"082082",
   56912 => x"082082",
   56913 => x"082082",
   56914 => x"082082",
   56915 => x"082041",
   56916 => x"041041",
   56917 => x"041041",
   56918 => x"041041",
   56919 => x"041041",
   56920 => x"041041",
   56921 => x"041041",
   56922 => x"041041",
   56923 => x"041041",
   56924 => x"041041",
   56925 => x"041041",
   56926 => x"041041",
   56927 => x"041041",
   56928 => x"041041",
   56929 => x"041041",
   56930 => x"041041",
   56931 => x"041041",
   56932 => x"041041",
   56933 => x"041041",
   56934 => x"041041",
   56935 => x"041041",
   56936 => x"041041",
   56937 => x"041041",
   56938 => x"041000",
   56939 => x"000000",
   56940 => x"000000",
   56941 => x"000000",
   56942 => x"000000",
   56943 => x"000000",
   56944 => x"000000",
   56945 => x"000000",
   56946 => x"000000",
   56947 => x"000000",
   56948 => x"000000",
   56949 => x"00057f",
   56950 => x"ffffff",
   56951 => x"ffffff",
   56952 => x"ffffff",
   56953 => x"ffffff",
   56954 => x"ffffff",
   56955 => x"ffffff",
   56956 => x"ffffff",
   56957 => x"ffffff",
   56958 => x"ffffff",
   56959 => x"ffffff",
   56960 => x"ffffff",
   56961 => x"ffffff",
   56962 => x"ffffff",
   56963 => x"ffffff",
   56964 => x"ffffff",
   56965 => x"ffffff",
   56966 => x"ffffff",
   56967 => x"ffffff",
   56968 => x"ffffff",
   56969 => x"ffffff",
   56970 => x"ffffff",
   56971 => x"ffffff",
   56972 => x"ffffff",
   56973 => x"ffffff",
   56974 => x"ffffff",
   56975 => x"ffffff",
   56976 => x"ffffff",
   56977 => x"ffffff",
   56978 => x"ffffff",
   56979 => x"ffffff",
   56980 => x"ffffff",
   56981 => x"ffffff",
   56982 => x"ffffff",
   56983 => x"ffffff",
   56984 => x"ffffff",
   56985 => x"ffffff",
   56986 => x"ffffff",
   56987 => x"ffffff",
   56988 => x"ffffff",
   56989 => x"ffffff",
   56990 => x"ffffff",
   56991 => x"ffffff",
   56992 => x"ffffff",
   56993 => x"ffffff",
   56994 => x"ffffff",
   56995 => x"ffffff",
   56996 => x"ffffff",
   56997 => x"ffffff",
   56998 => x"ffffff",
   56999 => x"ffffff",
   57000 => x"ffffff",
   57001 => x"ffffff",
   57002 => x"ffffff",
   57003 => x"ffffff",
   57004 => x"ffffff",
   57005 => x"ffffff",
   57006 => x"ffffff",
   57007 => x"ffffff",
   57008 => x"ffffff",
   57009 => x"ffffff",
   57010 => x"ffffff",
   57011 => x"ffffff",
   57012 => x"ffffff",
   57013 => x"ffffff",
   57014 => x"ffffff",
   57015 => x"ffffff",
   57016 => x"ffffff",
   57017 => x"ffffff",
   57018 => x"ffffff",
   57019 => x"ffffff",
   57020 => x"ffffff",
   57021 => x"ffffff",
   57022 => x"ffffff",
   57023 => x"ffffff",
   57024 => x"ffffff",
   57025 => x"ffffff",
   57026 => x"ffffff",
   57027 => x"ffffff",
   57028 => x"ffffff",
   57029 => x"fffa95",
   57030 => x"abffff",
   57031 => x"ffffff",
   57032 => x"ffffff",
   57033 => x"ffffff",
   57034 => x"ffffff",
   57035 => x"ffffff",
   57036 => x"ffffff",
   57037 => x"ffffff",
   57038 => x"ffffff",
   57039 => x"ffffff",
   57040 => x"ffffff",
   57041 => x"fffac3",
   57042 => x"0c30c3",
   57043 => x"0c30c3",
   57044 => x"0c30c3",
   57045 => x"0c30c3",
   57046 => x"0c30c3",
   57047 => x"0c30c3",
   57048 => x"0c30c3",
   57049 => x"0c30c3",
   57050 => x"0c30c3",
   57051 => x"0c30c3",
   57052 => x"0c30c3",
   57053 => x"082082",
   57054 => x"082082",
   57055 => x"082082",
   57056 => x"082082",
   57057 => x"082082",
   57058 => x"082082",
   57059 => x"082082",
   57060 => x"082082",
   57061 => x"082082",
   57062 => x"082082",
   57063 => x"082082",
   57064 => x"082082",
   57065 => x"082082",
   57066 => x"082082",
   57067 => x"082082",
   57068 => x"082082",
   57069 => x"082082",
   57070 => x"082082",
   57071 => x"082082",
   57072 => x"082082",
   57073 => x"082082",
   57074 => x"082082",
   57075 => x"082041",
   57076 => x"041041",
   57077 => x"041041",
   57078 => x"041041",
   57079 => x"041041",
   57080 => x"041041",
   57081 => x"041041",
   57082 => x"041041",
   57083 => x"041041",
   57084 => x"041041",
   57085 => x"041041",
   57086 => x"041041",
   57087 => x"041041",
   57088 => x"041041",
   57089 => x"041041",
   57090 => x"041041",
   57091 => x"041041",
   57092 => x"041041",
   57093 => x"041041",
   57094 => x"041041",
   57095 => x"041041",
   57096 => x"041041",
   57097 => x"041041",
   57098 => x"041000",
   57099 => x"000000",
   57100 => x"000000",
   57101 => x"000000",
   57102 => x"000000",
   57103 => x"000000",
   57104 => x"000000",
   57105 => x"000000",
   57106 => x"000000",
   57107 => x"000000",
   57108 => x"000000",
   57109 => x"00057f",
   57110 => x"ffffff",
   57111 => x"ffffff",
   57112 => x"ffffff",
   57113 => x"ffffff",
   57114 => x"ffffff",
   57115 => x"ffffff",
   57116 => x"ffffff",
   57117 => x"ffffff",
   57118 => x"ffffff",
   57119 => x"ffffff",
   57120 => x"ffffff",
   57121 => x"ffffff",
   57122 => x"ffffff",
   57123 => x"ffffff",
   57124 => x"ffffff",
   57125 => x"ffffff",
   57126 => x"ffffff",
   57127 => x"ffffff",
   57128 => x"ffffff",
   57129 => x"ffffff",
   57130 => x"ffffff",
   57131 => x"ffffff",
   57132 => x"ffffff",
   57133 => x"ffffff",
   57134 => x"ffffff",
   57135 => x"ffffff",
   57136 => x"ffffff",
   57137 => x"ffffff",
   57138 => x"ffffff",
   57139 => x"ffffff",
   57140 => x"ffffff",
   57141 => x"ffffff",
   57142 => x"ffffff",
   57143 => x"ffffff",
   57144 => x"ffffff",
   57145 => x"ffffff",
   57146 => x"ffffff",
   57147 => x"ffffff",
   57148 => x"ffffff",
   57149 => x"ffffff",
   57150 => x"ffffff",
   57151 => x"ffffff",
   57152 => x"ffffff",
   57153 => x"ffffff",
   57154 => x"ffffff",
   57155 => x"ffffff",
   57156 => x"ffffff",
   57157 => x"ffffff",
   57158 => x"ffffff",
   57159 => x"ffffff",
   57160 => x"ffffff",
   57161 => x"ffffff",
   57162 => x"ffffff",
   57163 => x"ffffff",
   57164 => x"ffffff",
   57165 => x"ffffff",
   57166 => x"ffffff",
   57167 => x"ffffff",
   57168 => x"ffffff",
   57169 => x"ffffff",
   57170 => x"ffffff",
   57171 => x"ffffff",
   57172 => x"ffffff",
   57173 => x"ffffff",
   57174 => x"ffffff",
   57175 => x"ffffff",
   57176 => x"ffffff",
   57177 => x"ffffff",
   57178 => x"ffffff",
   57179 => x"ffffff",
   57180 => x"ffffff",
   57181 => x"ffffff",
   57182 => x"ffffff",
   57183 => x"ffffff",
   57184 => x"ffffff",
   57185 => x"ffffff",
   57186 => x"ffffff",
   57187 => x"ffffff",
   57188 => x"ffffff",
   57189 => x"fffa95",
   57190 => x"abffff",
   57191 => x"ffffff",
   57192 => x"ffffff",
   57193 => x"ffffff",
   57194 => x"ffffff",
   57195 => x"ffffff",
   57196 => x"ffffff",
   57197 => x"ffffff",
   57198 => x"ffffff",
   57199 => x"ffffff",
   57200 => x"ffffff",
   57201 => x"fffac3",
   57202 => x"0c30c3",
   57203 => x"0c30c3",
   57204 => x"0c30c3",
   57205 => x"0c30c3",
   57206 => x"0c30c3",
   57207 => x"0c30c3",
   57208 => x"0c30c3",
   57209 => x"0c30c3",
   57210 => x"0c30c3",
   57211 => x"0c30c3",
   57212 => x"0c30c3",
   57213 => x"082082",
   57214 => x"082082",
   57215 => x"082082",
   57216 => x"082082",
   57217 => x"082082",
   57218 => x"082082",
   57219 => x"082082",
   57220 => x"082082",
   57221 => x"082082",
   57222 => x"082082",
   57223 => x"082082",
   57224 => x"082082",
   57225 => x"082082",
   57226 => x"082082",
   57227 => x"082082",
   57228 => x"082082",
   57229 => x"082082",
   57230 => x"082082",
   57231 => x"082082",
   57232 => x"082082",
   57233 => x"082082",
   57234 => x"082082",
   57235 => x"082041",
   57236 => x"041041",
   57237 => x"041041",
   57238 => x"041041",
   57239 => x"041041",
   57240 => x"041041",
   57241 => x"041041",
   57242 => x"041041",
   57243 => x"041041",
   57244 => x"041041",
   57245 => x"041041",
   57246 => x"041041",
   57247 => x"041041",
   57248 => x"041041",
   57249 => x"041041",
   57250 => x"041041",
   57251 => x"041041",
   57252 => x"041041",
   57253 => x"041041",
   57254 => x"041041",
   57255 => x"041041",
   57256 => x"041041",
   57257 => x"041041",
   57258 => x"041000",
   57259 => x"000000",
   57260 => x"000000",
   57261 => x"000000",
   57262 => x"000000",
   57263 => x"000000",
   57264 => x"000000",
   57265 => x"000000",
   57266 => x"000000",
   57267 => x"000000",
   57268 => x"000000",
   57269 => x"00057f",
   57270 => x"ffffff",
   57271 => x"ffffff",
   57272 => x"ffffff",
   57273 => x"ffffff",
   57274 => x"ffffff",
   57275 => x"ffffff",
   57276 => x"ffffff",
   57277 => x"ffffff",
   57278 => x"ffffff",
   57279 => x"ffffff",
   57280 => x"ffffff",
   57281 => x"ffffff",
   57282 => x"ffffff",
   57283 => x"ffffff",
   57284 => x"ffffff",
   57285 => x"ffffff",
   57286 => x"ffffff",
   57287 => x"ffffff",
   57288 => x"ffffff",
   57289 => x"ffffff",
   57290 => x"ffffff",
   57291 => x"ffffff",
   57292 => x"ffffff",
   57293 => x"ffffff",
   57294 => x"ffffff",
   57295 => x"ffffff",
   57296 => x"ffffff",
   57297 => x"ffffff",
   57298 => x"ffffff",
   57299 => x"ffffff",
   57300 => x"ffffff",
   57301 => x"ffffff",
   57302 => x"ffffff",
   57303 => x"ffffff",
   57304 => x"ffffff",
   57305 => x"ffffff",
   57306 => x"ffffff",
   57307 => x"ffffff",
   57308 => x"ffffff",
   57309 => x"ffffff",
   57310 => x"ffffff",
   57311 => x"ffffff",
   57312 => x"ffffff",
   57313 => x"ffffff",
   57314 => x"ffffff",
   57315 => x"ffffff",
   57316 => x"ffffff",
   57317 => x"ffffff",
   57318 => x"ffffff",
   57319 => x"ffffff",
   57320 => x"ffffff",
   57321 => x"ffffff",
   57322 => x"ffffff",
   57323 => x"ffffff",
   57324 => x"ffffff",
   57325 => x"ffffff",
   57326 => x"ffffff",
   57327 => x"ffffff",
   57328 => x"ffffff",
   57329 => x"ffffff",
   57330 => x"ffffff",
   57331 => x"ffffff",
   57332 => x"ffffff",
   57333 => x"ffffff",
   57334 => x"ffffff",
   57335 => x"ffffff",
   57336 => x"ffffff",
   57337 => x"ffffff",
   57338 => x"ffffff",
   57339 => x"ffffff",
   57340 => x"ffffff",
   57341 => x"ffffff",
   57342 => x"ffffff",
   57343 => x"ffffff",
   57344 => x"ffffff",
   57345 => x"ffffff",
   57346 => x"ffffff",
   57347 => x"ffffff",
   57348 => x"ffffff",
   57349 => x"fffa95",
   57350 => x"abffff",
   57351 => x"ffffff",
   57352 => x"ffffff",
   57353 => x"ffffff",
   57354 => x"ffffff",
   57355 => x"ffffff",
   57356 => x"ffffff",
   57357 => x"ffffff",
   57358 => x"ffffff",
   57359 => x"ffffff",
   57360 => x"ffffff",
   57361 => x"fffac3",
   57362 => x"0c30c3",
   57363 => x"0c30c3",
   57364 => x"0c30c3",
   57365 => x"0c30c3",
   57366 => x"0c30c3",
   57367 => x"0c30c3",
   57368 => x"0c30c3",
   57369 => x"0c30c3",
   57370 => x"0c30c3",
   57371 => x"0c30c3",
   57372 => x"0c30c3",
   57373 => x"082082",
   57374 => x"082082",
   57375 => x"082082",
   57376 => x"082082",
   57377 => x"082082",
   57378 => x"082082",
   57379 => x"082082",
   57380 => x"082082",
   57381 => x"082082",
   57382 => x"082082",
   57383 => x"082082",
   57384 => x"082082",
   57385 => x"082082",
   57386 => x"082082",
   57387 => x"082082",
   57388 => x"082082",
   57389 => x"082082",
   57390 => x"082082",
   57391 => x"082082",
   57392 => x"082082",
   57393 => x"082082",
   57394 => x"082082",
   57395 => x"082041",
   57396 => x"041041",
   57397 => x"041041",
   57398 => x"041041",
   57399 => x"041041",
   57400 => x"041041",
   57401 => x"041041",
   57402 => x"041041",
   57403 => x"041041",
   57404 => x"041041",
   57405 => x"041041",
   57406 => x"041041",
   57407 => x"041041",
   57408 => x"041041",
   57409 => x"041041",
   57410 => x"041041",
   57411 => x"041041",
   57412 => x"041041",
   57413 => x"041041",
   57414 => x"041041",
   57415 => x"041041",
   57416 => x"041041",
   57417 => x"041041",
   57418 => x"041000",
   57419 => x"000000",
   57420 => x"000000",
   57421 => x"000000",
   57422 => x"000000",
   57423 => x"000000",
   57424 => x"000000",
   57425 => x"000000",
   57426 => x"000000",
   57427 => x"000000",
   57428 => x"000000",
   57429 => x"00057f",
   57430 => x"ffffff",
   57431 => x"ffffff",
   57432 => x"ffffff",
   57433 => x"ffffff",
   57434 => x"ffffff",
   57435 => x"ffffff",
   57436 => x"ffffff",
   57437 => x"ffffff",
   57438 => x"ffffff",
   57439 => x"ffffff",
   57440 => x"ffffff",
   57441 => x"ffffff",
   57442 => x"ffffff",
   57443 => x"ffffff",
   57444 => x"ffffff",
   57445 => x"ffffff",
   57446 => x"ffffff",
   57447 => x"ffffff",
   57448 => x"ffffff",
   57449 => x"ffffff",
   57450 => x"ffffff",
   57451 => x"ffffff",
   57452 => x"ffffff",
   57453 => x"ffffff",
   57454 => x"ffffff",
   57455 => x"ffffff",
   57456 => x"ffffff",
   57457 => x"ffffff",
   57458 => x"ffffff",
   57459 => x"ffffff",
   57460 => x"ffffff",
   57461 => x"ffffff",
   57462 => x"ffffff",
   57463 => x"ffffff",
   57464 => x"ffffff",
   57465 => x"ffffff",
   57466 => x"ffffff",
   57467 => x"ffffff",
   57468 => x"ffffff",
   57469 => x"ffffff",
   57470 => x"ffffff",
   57471 => x"ffffff",
   57472 => x"ffffff",
   57473 => x"ffffff",
   57474 => x"ffffff",
   57475 => x"ffffff",
   57476 => x"ffffff",
   57477 => x"ffffff",
   57478 => x"ffffff",
   57479 => x"ffffff",
   57480 => x"ffffff",
   57481 => x"ffffff",
   57482 => x"ffffff",
   57483 => x"ffffff",
   57484 => x"ffffff",
   57485 => x"ffffff",
   57486 => x"ffffff",
   57487 => x"ffffff",
   57488 => x"ffffff",
   57489 => x"ffffff",
   57490 => x"ffffff",
   57491 => x"ffffff",
   57492 => x"ffffff",
   57493 => x"ffffff",
   57494 => x"ffffff",
   57495 => x"ffffff",
   57496 => x"ffffff",
   57497 => x"ffffff",
   57498 => x"ffffff",
   57499 => x"ffffff",
   57500 => x"ffffff",
   57501 => x"ffffff",
   57502 => x"ffffff",
   57503 => x"ffffff",
   57504 => x"ffffff",
   57505 => x"ffffff",
   57506 => x"ffffff",
   57507 => x"ffffff",
   57508 => x"ffffff",
   57509 => x"fffa95",
   57510 => x"abffff",
   57511 => x"ffffff",
   57512 => x"ffffff",
   57513 => x"ffffff",
   57514 => x"ffffff",
   57515 => x"ffffff",
   57516 => x"ffffff",
   57517 => x"ffffff",
   57518 => x"ffffff",
   57519 => x"ffffff",
   57520 => x"ffffff",
   57521 => x"fffac3",
   57522 => x"0c30c3",
   57523 => x"0c30c3",
   57524 => x"0c30c3",
   57525 => x"0c30c3",
   57526 => x"0c30c3",
   57527 => x"0c30c3",
   57528 => x"0c30c3",
   57529 => x"0c30c3",
   57530 => x"0c30c3",
   57531 => x"0c30c3",
   57532 => x"0c30c3",
   57533 => x"082082",
   57534 => x"082082",
   57535 => x"082082",
   57536 => x"082082",
   57537 => x"082082",
   57538 => x"082082",
   57539 => x"082082",
   57540 => x"082082",
   57541 => x"082082",
   57542 => x"082082",
   57543 => x"082082",
   57544 => x"082082",
   57545 => x"082082",
   57546 => x"082082",
   57547 => x"082082",
   57548 => x"082082",
   57549 => x"082082",
   57550 => x"082082",
   57551 => x"082082",
   57552 => x"082082",
   57553 => x"082082",
   57554 => x"082082",
   57555 => x"082041",
   57556 => x"041041",
   57557 => x"041041",
   57558 => x"041041",
   57559 => x"041041",
   57560 => x"041041",
   57561 => x"041041",
   57562 => x"041041",
   57563 => x"041041",
   57564 => x"041041",
   57565 => x"041041",
   57566 => x"041041",
   57567 => x"041041",
   57568 => x"041041",
   57569 => x"041041",
   57570 => x"041041",
   57571 => x"041041",
   57572 => x"041041",
   57573 => x"041041",
   57574 => x"041041",
   57575 => x"041041",
   57576 => x"041041",
   57577 => x"041041",
   57578 => x"041000",
   57579 => x"000000",
   57580 => x"000000",
   57581 => x"000000",
   57582 => x"000000",
   57583 => x"000000",
   57584 => x"000000",
   57585 => x"000000",
   57586 => x"000000",
   57587 => x"000000",
   57588 => x"000000",
   57589 => x"00057f",
   57590 => x"ffffff",
   57591 => x"ffffff",
   57592 => x"ffffff",
   57593 => x"ffffff",
   57594 => x"ffffff",
   57595 => x"ffffff",
   57596 => x"ffffff",
   57597 => x"ffffff",
   57598 => x"ffffff",
   57599 => x"ffffff",
   57600 => x"ffffff",
   57601 => x"ffffff",
   57602 => x"ffffff",
   57603 => x"ffffff",
   57604 => x"ffffff",
   57605 => x"ffffff",
   57606 => x"ffffff",
   57607 => x"ffffff",
   57608 => x"ffffff",
   57609 => x"ffffff",
   57610 => x"ffffff",
   57611 => x"ffffff",
   57612 => x"ffffff",
   57613 => x"ffffff",
   57614 => x"ffffff",
   57615 => x"ffffff",
   57616 => x"ffffff",
   57617 => x"ffffff",
   57618 => x"ffffff",
   57619 => x"ffffff",
   57620 => x"ffffff",
   57621 => x"ffffff",
   57622 => x"ffffff",
   57623 => x"ffffff",
   57624 => x"ffffff",
   57625 => x"ffffff",
   57626 => x"ffffff",
   57627 => x"ffffff",
   57628 => x"ffffff",
   57629 => x"ffffff",
   57630 => x"ffffff",
   57631 => x"ffffff",
   57632 => x"ffffff",
   57633 => x"ffffff",
   57634 => x"ffffff",
   57635 => x"ffffff",
   57636 => x"ffffff",
   57637 => x"ffffff",
   57638 => x"ffffff",
   57639 => x"ffffff",
   57640 => x"ffffff",
   57641 => x"ffffff",
   57642 => x"ffffff",
   57643 => x"ffffff",
   57644 => x"ffffff",
   57645 => x"ffffff",
   57646 => x"ffffff",
   57647 => x"ffffff",
   57648 => x"ffffff",
   57649 => x"ffffff",
   57650 => x"ffffff",
   57651 => x"ffffff",
   57652 => x"ffffff",
   57653 => x"ffffff",
   57654 => x"ffffff",
   57655 => x"ffffff",
   57656 => x"ffffff",
   57657 => x"ffffff",
   57658 => x"ffffff",
   57659 => x"ffffff",
   57660 => x"ffffff",
   57661 => x"ffffff",
   57662 => x"ffffff",
   57663 => x"ffffff",
   57664 => x"ffffff",
   57665 => x"ffffff",
   57666 => x"ffffff",
   57667 => x"ffffff",
   57668 => x"ffffff",
   57669 => x"fffa95",
   57670 => x"abffff",
   57671 => x"ffffff",
   57672 => x"ffffff",
   57673 => x"ffffff",
   57674 => x"ffffff",
   57675 => x"ffffff",
   57676 => x"ffffff",
   57677 => x"ffffff",
   57678 => x"ffffff",
   57679 => x"ffffff",
   57680 => x"ffffff",
   57681 => x"fffac3",
   57682 => x"0c30c3",
   57683 => x"0c30c3",
   57684 => x"0c30c3",
   57685 => x"0c30c3",
   57686 => x"0c30c3",
   57687 => x"0c30c3",
   57688 => x"0c30c3",
   57689 => x"0c30c3",
   57690 => x"0c30c3",
   57691 => x"0c30c3",
   57692 => x"0c30c3",
   57693 => x"082082",
   57694 => x"082082",
   57695 => x"082082",
   57696 => x"082082",
   57697 => x"082082",
   57698 => x"082082",
   57699 => x"082082",
   57700 => x"082082",
   57701 => x"082082",
   57702 => x"082082",
   57703 => x"082082",
   57704 => x"082082",
   57705 => x"082082",
   57706 => x"082082",
   57707 => x"082082",
   57708 => x"082082",
   57709 => x"082082",
   57710 => x"082082",
   57711 => x"082082",
   57712 => x"082082",
   57713 => x"082082",
   57714 => x"082082",
   57715 => x"082041",
   57716 => x"041041",
   57717 => x"041041",
   57718 => x"041041",
   57719 => x"041041",
   57720 => x"041041",
   57721 => x"041041",
   57722 => x"041041",
   57723 => x"041041",
   57724 => x"041041",
   57725 => x"041041",
   57726 => x"041041",
   57727 => x"041041",
   57728 => x"041041",
   57729 => x"041041",
   57730 => x"041041",
   57731 => x"041041",
   57732 => x"041041",
   57733 => x"041041",
   57734 => x"041041",
   57735 => x"041041",
   57736 => x"041041",
   57737 => x"041041",
   57738 => x"041000",
   57739 => x"000000",
   57740 => x"000000",
   57741 => x"000000",
   57742 => x"000000",
   57743 => x"000000",
   57744 => x"000000",
   57745 => x"000000",
   57746 => x"000000",
   57747 => x"000000",
   57748 => x"000000",
   57749 => x"00057f",
   57750 => x"ffffff",
   57751 => x"ffffff",
   57752 => x"ffffff",
   57753 => x"ffffff",
   57754 => x"ffffff",
   57755 => x"ffffff",
   57756 => x"ffffff",
   57757 => x"ffffff",
   57758 => x"ffffff",
   57759 => x"ffffff",
   57760 => x"ffffff",
   57761 => x"ffffff",
   57762 => x"ffffff",
   57763 => x"ffffff",
   57764 => x"ffffff",
   57765 => x"ffffff",
   57766 => x"ffffff",
   57767 => x"ffffff",
   57768 => x"ffffff",
   57769 => x"ffffff",
   57770 => x"ffffff",
   57771 => x"ffffff",
   57772 => x"ffffff",
   57773 => x"ffffff",
   57774 => x"ffffff",
   57775 => x"ffffff",
   57776 => x"ffffff",
   57777 => x"ffffff",
   57778 => x"ffffff",
   57779 => x"ffffff",
   57780 => x"ffffff",
   57781 => x"ffffff",
   57782 => x"ffffff",
   57783 => x"ffffff",
   57784 => x"ffffff",
   57785 => x"ffffff",
   57786 => x"ffffff",
   57787 => x"ffffff",
   57788 => x"ffffff",
   57789 => x"ffffff",
   57790 => x"ffffff",
   57791 => x"ffffff",
   57792 => x"ffffff",
   57793 => x"ffffff",
   57794 => x"ffffff",
   57795 => x"ffffff",
   57796 => x"ffffff",
   57797 => x"ffffff",
   57798 => x"ffffff",
   57799 => x"ffffff",
   57800 => x"ffffff",
   57801 => x"ffffff",
   57802 => x"ffffff",
   57803 => x"ffffff",
   57804 => x"ffffff",
   57805 => x"ffffff",
   57806 => x"ffffff",
   57807 => x"ffffff",
   57808 => x"ffffff",
   57809 => x"ffffff",
   57810 => x"ffffff",
   57811 => x"ffffff",
   57812 => x"ffffff",
   57813 => x"ffffff",
   57814 => x"ffffff",
   57815 => x"ffffff",
   57816 => x"ffffff",
   57817 => x"ffffff",
   57818 => x"ffffff",
   57819 => x"ffffff",
   57820 => x"ffffff",
   57821 => x"ffffff",
   57822 => x"ffffff",
   57823 => x"ffffff",
   57824 => x"ffffff",
   57825 => x"ffffff",
   57826 => x"ffffff",
   57827 => x"ffffff",
   57828 => x"ffffff",
   57829 => x"fffa95",
   57830 => x"abffff",
   57831 => x"ffffff",
   57832 => x"ffffff",
   57833 => x"ffffff",
   57834 => x"ffffff",
   57835 => x"ffffff",
   57836 => x"ffffff",
   57837 => x"ffffff",
   57838 => x"ffffff",
   57839 => x"ffffff",
   57840 => x"ffffff",
   57841 => x"fffac3",
   57842 => x"0c30c3",
   57843 => x"0c30c3",
   57844 => x"0c30c3",
   57845 => x"0c30c3",
   57846 => x"0c30c3",
   57847 => x"0c30c3",
   57848 => x"0c30c3",
   57849 => x"0c30c3",
   57850 => x"0c30c3",
   57851 => x"0c30c3",
   57852 => x"0c30c3",
   57853 => x"082082",
   57854 => x"082082",
   57855 => x"082082",
   57856 => x"082082",
   57857 => x"082082",
   57858 => x"082082",
   57859 => x"082082",
   57860 => x"082082",
   57861 => x"082082",
   57862 => x"082082",
   57863 => x"082082",
   57864 => x"082082",
   57865 => x"082082",
   57866 => x"082082",
   57867 => x"082082",
   57868 => x"082082",
   57869 => x"082082",
   57870 => x"082082",
   57871 => x"082082",
   57872 => x"082082",
   57873 => x"082082",
   57874 => x"082082",
   57875 => x"082041",
   57876 => x"041041",
   57877 => x"041041",
   57878 => x"041041",
   57879 => x"041041",
   57880 => x"041041",
   57881 => x"041041",
   57882 => x"041041",
   57883 => x"041041",
   57884 => x"041041",
   57885 => x"041041",
   57886 => x"041041",
   57887 => x"041041",
   57888 => x"041041",
   57889 => x"041041",
   57890 => x"041041",
   57891 => x"041041",
   57892 => x"041041",
   57893 => x"041041",
   57894 => x"041041",
   57895 => x"041041",
   57896 => x"041041",
   57897 => x"041041",
   57898 => x"041000",
   57899 => x"000000",
   57900 => x"000000",
   57901 => x"000000",
   57902 => x"000000",
   57903 => x"000000",
   57904 => x"000000",
   57905 => x"000000",
   57906 => x"000000",
   57907 => x"000000",
   57908 => x"000000",
   57909 => x"00057f",
   57910 => x"ffffff",
   57911 => x"ffffff",
   57912 => x"ffffff",
   57913 => x"ffffff",
   57914 => x"ffffff",
   57915 => x"ffffff",
   57916 => x"ffffff",
   57917 => x"ffffff",
   57918 => x"ffffff",
   57919 => x"ffffff",
   57920 => x"ffffff",
   57921 => x"ffffff",
   57922 => x"ffffff",
   57923 => x"ffffff",
   57924 => x"ffffff",
   57925 => x"ffffff",
   57926 => x"ffffff",
   57927 => x"ffffff",
   57928 => x"ffffff",
   57929 => x"ffffff",
   57930 => x"ffffff",
   57931 => x"ffffff",
   57932 => x"ffffff",
   57933 => x"ffffff",
   57934 => x"ffffff",
   57935 => x"ffffff",
   57936 => x"ffffff",
   57937 => x"ffffff",
   57938 => x"ffffff",
   57939 => x"ffffff",
   57940 => x"ffffff",
   57941 => x"ffffff",
   57942 => x"ffffff",
   57943 => x"ffffff",
   57944 => x"ffffff",
   57945 => x"ffffff",
   57946 => x"ffffff",
   57947 => x"ffffff",
   57948 => x"ffffff",
   57949 => x"ffffff",
   57950 => x"ffffff",
   57951 => x"ffffff",
   57952 => x"ffffff",
   57953 => x"ffffff",
   57954 => x"ffffff",
   57955 => x"ffffff",
   57956 => x"ffffff",
   57957 => x"ffffff",
   57958 => x"ffffff",
   57959 => x"ffffff",
   57960 => x"ffffff",
   57961 => x"ffffff",
   57962 => x"ffffff",
   57963 => x"ffffff",
   57964 => x"ffffff",
   57965 => x"ffffff",
   57966 => x"ffffff",
   57967 => x"ffffff",
   57968 => x"ffffff",
   57969 => x"ffffff",
   57970 => x"ffffff",
   57971 => x"ffffff",
   57972 => x"ffffff",
   57973 => x"ffffff",
   57974 => x"ffffff",
   57975 => x"ffffff",
   57976 => x"ffffff",
   57977 => x"ffffff",
   57978 => x"ffffff",
   57979 => x"ffffff",
   57980 => x"ffffff",
   57981 => x"ffffff",
   57982 => x"ffffff",
   57983 => x"ffffff",
   57984 => x"ffffff",
   57985 => x"ffffff",
   57986 => x"ffffff",
   57987 => x"ffffff",
   57988 => x"ffffff",
   57989 => x"fffa95",
   57990 => x"abffff",
   57991 => x"ffffff",
   57992 => x"ffffff",
   57993 => x"ffffff",
   57994 => x"ffffff",
   57995 => x"ffffff",
   57996 => x"ffffff",
   57997 => x"ffffff",
   57998 => x"ffffff",
   57999 => x"ffffff",
   58000 => x"ffffff",
   58001 => x"fffac3",
   58002 => x"0c30c3",
   58003 => x"0c30c3",
   58004 => x"0c30c3",
   58005 => x"0c30c3",
   58006 => x"0c30c3",
   58007 => x"0c30c3",
   58008 => x"0c30c3",
   58009 => x"0c30c3",
   58010 => x"0c30c3",
   58011 => x"0c30c3",
   58012 => x"0c30c3",
   58013 => x"082082",
   58014 => x"082082",
   58015 => x"082082",
   58016 => x"082082",
   58017 => x"082082",
   58018 => x"082082",
   58019 => x"082082",
   58020 => x"082082",
   58021 => x"082082",
   58022 => x"082082",
   58023 => x"082082",
   58024 => x"082082",
   58025 => x"082082",
   58026 => x"082082",
   58027 => x"082082",
   58028 => x"082082",
   58029 => x"082082",
   58030 => x"082082",
   58031 => x"082082",
   58032 => x"082082",
   58033 => x"082082",
   58034 => x"082082",
   58035 => x"082041",
   58036 => x"041041",
   58037 => x"041041",
   58038 => x"041041",
   58039 => x"041041",
   58040 => x"041041",
   58041 => x"041041",
   58042 => x"041041",
   58043 => x"041041",
   58044 => x"041041",
   58045 => x"041041",
   58046 => x"041041",
   58047 => x"041041",
   58048 => x"041041",
   58049 => x"041041",
   58050 => x"041041",
   58051 => x"041041",
   58052 => x"041041",
   58053 => x"041041",
   58054 => x"041041",
   58055 => x"041041",
   58056 => x"041041",
   58057 => x"041041",
   58058 => x"041000",
   58059 => x"000000",
   58060 => x"000000",
   58061 => x"000000",
   58062 => x"000000",
   58063 => x"000000",
   58064 => x"000000",
   58065 => x"000000",
   58066 => x"000000",
   58067 => x"000000",
   58068 => x"000000",
   58069 => x"00057f",
   58070 => x"ffffff",
   58071 => x"ffffff",
   58072 => x"ffffff",
   58073 => x"ffffff",
   58074 => x"ffffff",
   58075 => x"ffffff",
   58076 => x"ffffff",
   58077 => x"ffffff",
   58078 => x"ffffff",
   58079 => x"ffffff",
   58080 => x"ffffff",
   58081 => x"ffffff",
   58082 => x"ffffff",
   58083 => x"ffffff",
   58084 => x"ffffff",
   58085 => x"ffffff",
   58086 => x"ffffff",
   58087 => x"ffffff",
   58088 => x"ffffff",
   58089 => x"ffffff",
   58090 => x"ffffff",
   58091 => x"ffffff",
   58092 => x"ffffff",
   58093 => x"ffffff",
   58094 => x"ffffff",
   58095 => x"ffffff",
   58096 => x"ffffff",
   58097 => x"ffffff",
   58098 => x"ffffff",
   58099 => x"ffffff",
   58100 => x"ffffff",
   58101 => x"ffffff",
   58102 => x"ffffff",
   58103 => x"ffffff",
   58104 => x"ffffff",
   58105 => x"ffffff",
   58106 => x"ffffff",
   58107 => x"ffffff",
   58108 => x"ffffff",
   58109 => x"ffffff",
   58110 => x"ffffff",
   58111 => x"ffffff",
   58112 => x"ffffff",
   58113 => x"ffffff",
   58114 => x"ffffff",
   58115 => x"ffffff",
   58116 => x"ffffff",
   58117 => x"ffffff",
   58118 => x"ffffff",
   58119 => x"ffffff",
   58120 => x"ffffff",
   58121 => x"ffffff",
   58122 => x"ffffff",
   58123 => x"ffffff",
   58124 => x"ffffff",
   58125 => x"ffffff",
   58126 => x"ffffff",
   58127 => x"ffffff",
   58128 => x"ffffff",
   58129 => x"ffffff",
   58130 => x"ffffff",
   58131 => x"ffffff",
   58132 => x"ffffff",
   58133 => x"ffffff",
   58134 => x"ffffff",
   58135 => x"ffffff",
   58136 => x"ffffff",
   58137 => x"ffffff",
   58138 => x"ffffff",
   58139 => x"ffffff",
   58140 => x"ffffff",
   58141 => x"ffffff",
   58142 => x"ffffff",
   58143 => x"ffffff",
   58144 => x"ffffff",
   58145 => x"ffffff",
   58146 => x"ffffff",
   58147 => x"ffffff",
   58148 => x"ffffff",
   58149 => x"fffa95",
   58150 => x"abffff",
   58151 => x"ffffff",
   58152 => x"ffffff",
   58153 => x"ffffff",
   58154 => x"ffffff",
   58155 => x"ffffff",
   58156 => x"ffffff",
   58157 => x"ffffff",
   58158 => x"ffffff",
   58159 => x"ffffff",
   58160 => x"ffffff",
   58161 => x"fffac3",
   58162 => x"0c30c3",
   58163 => x"0c30c3",
   58164 => x"0c30c3",
   58165 => x"0c30c3",
   58166 => x"0c30c3",
   58167 => x"0c30c3",
   58168 => x"0c30c3",
   58169 => x"0c30c3",
   58170 => x"0c30c3",
   58171 => x"0c30c3",
   58172 => x"0c30c3",
   58173 => x"082082",
   58174 => x"082082",
   58175 => x"082082",
   58176 => x"082082",
   58177 => x"082082",
   58178 => x"082082",
   58179 => x"082082",
   58180 => x"082082",
   58181 => x"082082",
   58182 => x"082082",
   58183 => x"082082",
   58184 => x"082082",
   58185 => x"082082",
   58186 => x"082082",
   58187 => x"082082",
   58188 => x"082082",
   58189 => x"082082",
   58190 => x"082082",
   58191 => x"082082",
   58192 => x"082082",
   58193 => x"082082",
   58194 => x"082082",
   58195 => x"082041",
   58196 => x"041041",
   58197 => x"041041",
   58198 => x"041041",
   58199 => x"041041",
   58200 => x"041041",
   58201 => x"041041",
   58202 => x"041041",
   58203 => x"041041",
   58204 => x"041041",
   58205 => x"041041",
   58206 => x"041041",
   58207 => x"041041",
   58208 => x"041041",
   58209 => x"041041",
   58210 => x"041041",
   58211 => x"041041",
   58212 => x"041041",
   58213 => x"041041",
   58214 => x"041041",
   58215 => x"041041",
   58216 => x"041041",
   58217 => x"041041",
   58218 => x"041000",
   58219 => x"000000",
   58220 => x"000000",
   58221 => x"000000",
   58222 => x"000000",
   58223 => x"000000",
   58224 => x"000000",
   58225 => x"000000",
   58226 => x"000000",
   58227 => x"000000",
   58228 => x"000000",
   58229 => x"00057f",
   58230 => x"ffffff",
   58231 => x"ffffff",
   58232 => x"ffffff",
   58233 => x"ffffff",
   58234 => x"ffffff",
   58235 => x"ffffff",
   58236 => x"ffffff",
   58237 => x"ffffff",
   58238 => x"ffffff",
   58239 => x"ffffff",
   58240 => x"ffffff",
   58241 => x"ffffff",
   58242 => x"ffffff",
   58243 => x"ffffff",
   58244 => x"ffffff",
   58245 => x"ffffff",
   58246 => x"ffffff",
   58247 => x"ffffff",
   58248 => x"ffffff",
   58249 => x"ffffff",
   58250 => x"ffffff",
   58251 => x"ffffff",
   58252 => x"ffffff",
   58253 => x"ffffff",
   58254 => x"ffffff",
   58255 => x"ffffff",
   58256 => x"ffffff",
   58257 => x"ffffff",
   58258 => x"ffffff",
   58259 => x"ffffff",
   58260 => x"ffffff",
   58261 => x"ffffff",
   58262 => x"ffffff",
   58263 => x"ffffff",
   58264 => x"ffffff",
   58265 => x"ffffff",
   58266 => x"ffffff",
   58267 => x"ffffff",
   58268 => x"ffffff",
   58269 => x"ffffff",
   58270 => x"ffffff",
   58271 => x"ffffff",
   58272 => x"ffffff",
   58273 => x"ffffff",
   58274 => x"ffffff",
   58275 => x"ffffff",
   58276 => x"ffffff",
   58277 => x"ffffff",
   58278 => x"ffffff",
   58279 => x"ffffff",
   58280 => x"ffffff",
   58281 => x"ffffff",
   58282 => x"ffffff",
   58283 => x"ffffff",
   58284 => x"ffffff",
   58285 => x"ffffff",
   58286 => x"ffffff",
   58287 => x"ffffff",
   58288 => x"ffffff",
   58289 => x"ffffff",
   58290 => x"ffffff",
   58291 => x"ffffff",
   58292 => x"ffffff",
   58293 => x"ffffff",
   58294 => x"ffffff",
   58295 => x"ffffff",
   58296 => x"ffffff",
   58297 => x"ffffff",
   58298 => x"ffffff",
   58299 => x"ffffff",
   58300 => x"ffffff",
   58301 => x"ffffff",
   58302 => x"ffffff",
   58303 => x"ffffff",
   58304 => x"ffffff",
   58305 => x"ffffff",
   58306 => x"ffffff",
   58307 => x"ffffff",
   58308 => x"ffffff",
   58309 => x"fffa95",
   58310 => x"abffff",
   58311 => x"ffffff",
   58312 => x"ffffff",
   58313 => x"ffffff",
   58314 => x"ffffff",
   58315 => x"ffffff",
   58316 => x"ffffff",
   58317 => x"ffffff",
   58318 => x"ffffff",
   58319 => x"ffffff",
   58320 => x"ffffff",
   58321 => x"fffac3",
   58322 => x"0c30c3",
   58323 => x"0c30c3",
   58324 => x"0c30c3",
   58325 => x"0c30c3",
   58326 => x"0c30c3",
   58327 => x"0c30c3",
   58328 => x"0c30c3",
   58329 => x"0c30c3",
   58330 => x"0c30c3",
   58331 => x"0c30c3",
   58332 => x"0c30c3",
   58333 => x"082082",
   58334 => x"082082",
   58335 => x"082082",
   58336 => x"082082",
   58337 => x"082082",
   58338 => x"082082",
   58339 => x"082082",
   58340 => x"082082",
   58341 => x"082082",
   58342 => x"082082",
   58343 => x"082082",
   58344 => x"082082",
   58345 => x"082082",
   58346 => x"082082",
   58347 => x"082082",
   58348 => x"082082",
   58349 => x"082082",
   58350 => x"082082",
   58351 => x"082082",
   58352 => x"082082",
   58353 => x"082082",
   58354 => x"082082",
   58355 => x"082041",
   58356 => x"041041",
   58357 => x"041041",
   58358 => x"041041",
   58359 => x"041041",
   58360 => x"041041",
   58361 => x"041041",
   58362 => x"041041",
   58363 => x"041041",
   58364 => x"041041",
   58365 => x"041041",
   58366 => x"041041",
   58367 => x"041041",
   58368 => x"041041",
   58369 => x"041041",
   58370 => x"041041",
   58371 => x"041041",
   58372 => x"041041",
   58373 => x"041041",
   58374 => x"041041",
   58375 => x"041041",
   58376 => x"041041",
   58377 => x"041041",
   58378 => x"041000",
   58379 => x"000000",
   58380 => x"000000",
   58381 => x"000000",
   58382 => x"000000",
   58383 => x"000000",
   58384 => x"000000",
   58385 => x"000000",
   58386 => x"000000",
   58387 => x"000000",
   58388 => x"000000",
   58389 => x"00057f",
   58390 => x"ffffff",
   58391 => x"ffffff",
   58392 => x"ffffff",
   58393 => x"ffffff",
   58394 => x"ffffff",
   58395 => x"ffffff",
   58396 => x"ffffff",
   58397 => x"ffffff",
   58398 => x"ffffff",
   58399 => x"ffffff",
   58400 => x"ffffff",
   58401 => x"ffffff",
   58402 => x"ffffff",
   58403 => x"ffffff",
   58404 => x"ffffff",
   58405 => x"ffffff",
   58406 => x"ffffff",
   58407 => x"ffffff",
   58408 => x"ffffff",
   58409 => x"ffffff",
   58410 => x"ffffff",
   58411 => x"ffffff",
   58412 => x"ffffff",
   58413 => x"ffffff",
   58414 => x"ffffff",
   58415 => x"ffffff",
   58416 => x"ffffff",
   58417 => x"ffffff",
   58418 => x"ffffff",
   58419 => x"ffffff",
   58420 => x"ffffff",
   58421 => x"ffffff",
   58422 => x"ffffff",
   58423 => x"ffffff",
   58424 => x"ffffff",
   58425 => x"ffffff",
   58426 => x"ffffff",
   58427 => x"ffffff",
   58428 => x"ffffff",
   58429 => x"ffffff",
   58430 => x"ffffff",
   58431 => x"ffffff",
   58432 => x"ffffff",
   58433 => x"ffffff",
   58434 => x"ffffff",
   58435 => x"ffffff",
   58436 => x"ffffff",
   58437 => x"ffffff",
   58438 => x"ffffff",
   58439 => x"ffffff",
   58440 => x"ffffff",
   58441 => x"ffffff",
   58442 => x"ffffff",
   58443 => x"ffffff",
   58444 => x"ffffff",
   58445 => x"ffffff",
   58446 => x"ffffff",
   58447 => x"ffffff",
   58448 => x"ffffff",
   58449 => x"ffffff",
   58450 => x"ffffff",
   58451 => x"ffffff",
   58452 => x"ffffff",
   58453 => x"ffffff",
   58454 => x"ffffff",
   58455 => x"ffffff",
   58456 => x"ffffff",
   58457 => x"ffffff",
   58458 => x"ffffff",
   58459 => x"ffffff",
   58460 => x"ffffff",
   58461 => x"ffffff",
   58462 => x"ffffff",
   58463 => x"ffffff",
   58464 => x"ffffff",
   58465 => x"ffffff",
   58466 => x"ffffff",
   58467 => x"ffffff",
   58468 => x"ffffff",
   58469 => x"fffa95",
   58470 => x"abffff",
   58471 => x"ffffff",
   58472 => x"ffffff",
   58473 => x"ffffff",
   58474 => x"ffffff",
   58475 => x"ffffff",
   58476 => x"ffffff",
   58477 => x"ffffff",
   58478 => x"ffffff",
   58479 => x"ffffff",
   58480 => x"ffffff",
   58481 => x"fffac3",
   58482 => x"0c30c3",
   58483 => x"0c30c3",
   58484 => x"0c30c3",
   58485 => x"0c30c3",
   58486 => x"0c30c3",
   58487 => x"0c30c3",
   58488 => x"0c30c3",
   58489 => x"0c30c3",
   58490 => x"0c30c3",
   58491 => x"0c30c3",
   58492 => x"0c30c3",
   58493 => x"082082",
   58494 => x"082082",
   58495 => x"082082",
   58496 => x"082082",
   58497 => x"082082",
   58498 => x"082082",
   58499 => x"082082",
   58500 => x"082082",
   58501 => x"082082",
   58502 => x"082082",
   58503 => x"082082",
   58504 => x"082082",
   58505 => x"082082",
   58506 => x"082082",
   58507 => x"082082",
   58508 => x"082082",
   58509 => x"082082",
   58510 => x"082082",
   58511 => x"082082",
   58512 => x"082082",
   58513 => x"082082",
   58514 => x"082082",
   58515 => x"082041",
   58516 => x"041041",
   58517 => x"041041",
   58518 => x"041041",
   58519 => x"041041",
   58520 => x"041041",
   58521 => x"041041",
   58522 => x"041041",
   58523 => x"041041",
   58524 => x"041041",
   58525 => x"041041",
   58526 => x"041041",
   58527 => x"041041",
   58528 => x"041041",
   58529 => x"041041",
   58530 => x"041041",
   58531 => x"041041",
   58532 => x"041041",
   58533 => x"041041",
   58534 => x"041041",
   58535 => x"041041",
   58536 => x"041041",
   58537 => x"041041",
   58538 => x"041000",
   58539 => x"000000",
   58540 => x"000000",
   58541 => x"000000",
   58542 => x"000000",
   58543 => x"000000",
   58544 => x"000000",
   58545 => x"000000",
   58546 => x"000000",
   58547 => x"000000",
   58548 => x"000000",
   58549 => x"00057f",
   58550 => x"ffffff",
   58551 => x"ffffff",
   58552 => x"ffffff",
   58553 => x"ffffff",
   58554 => x"ffffff",
   58555 => x"ffffff",
   58556 => x"ffffff",
   58557 => x"ffffff",
   58558 => x"ffffff",
   58559 => x"ffffff",
   58560 => x"ffffff",
   58561 => x"ffffff",
   58562 => x"ffffff",
   58563 => x"ffffff",
   58564 => x"ffffff",
   58565 => x"ffffff",
   58566 => x"ffffff",
   58567 => x"ffffff",
   58568 => x"ffffff",
   58569 => x"ffffff",
   58570 => x"ffffff",
   58571 => x"ffffff",
   58572 => x"ffffff",
   58573 => x"ffffff",
   58574 => x"ffffff",
   58575 => x"ffffff",
   58576 => x"ffffff",
   58577 => x"ffffff",
   58578 => x"ffffff",
   58579 => x"ffffff",
   58580 => x"ffffff",
   58581 => x"ffffff",
   58582 => x"ffffff",
   58583 => x"ffffff",
   58584 => x"ffffff",
   58585 => x"ffffff",
   58586 => x"ffffff",
   58587 => x"ffffff",
   58588 => x"ffffff",
   58589 => x"ffffff",
   58590 => x"ffffff",
   58591 => x"ffffff",
   58592 => x"ffffff",
   58593 => x"ffffff",
   58594 => x"ffffff",
   58595 => x"ffffff",
   58596 => x"ffffff",
   58597 => x"ffffff",
   58598 => x"ffffff",
   58599 => x"ffffff",
   58600 => x"ffffff",
   58601 => x"ffffff",
   58602 => x"ffffff",
   58603 => x"ffffff",
   58604 => x"ffffff",
   58605 => x"ffffff",
   58606 => x"ffffff",
   58607 => x"ffffff",
   58608 => x"ffffff",
   58609 => x"ffffff",
   58610 => x"ffffff",
   58611 => x"ffffff",
   58612 => x"ffffff",
   58613 => x"ffffff",
   58614 => x"ffffff",
   58615 => x"ffffff",
   58616 => x"ffffff",
   58617 => x"ffffff",
   58618 => x"ffffff",
   58619 => x"ffffff",
   58620 => x"ffffff",
   58621 => x"ffffff",
   58622 => x"ffffff",
   58623 => x"ffffff",
   58624 => x"ffffff",
   58625 => x"ffffff",
   58626 => x"ffffff",
   58627 => x"ffffff",
   58628 => x"ffffff",
   58629 => x"fffa95",
   58630 => x"abffff",
   58631 => x"ffffff",
   58632 => x"ffffff",
   58633 => x"ffffff",
   58634 => x"ffffff",
   58635 => x"ffffff",
   58636 => x"ffffff",
   58637 => x"ffffff",
   58638 => x"ffffff",
   58639 => x"ffffff",
   58640 => x"ffffff",
   58641 => x"fffad7",
   58642 => x"0c30c3",
   58643 => x"0c30c3",
   58644 => x"0c30c3",
   58645 => x"0c30c3",
   58646 => x"0c30c3",
   58647 => x"0c30c3",
   58648 => x"0c30c3",
   58649 => x"0c30c3",
   58650 => x"0c30c3",
   58651 => x"0c30c3",
   58652 => x"0c30c3",
   58653 => x"0c30c3",
   58654 => x"082082",
   58655 => x"082082",
   58656 => x"082082",
   58657 => x"082082",
   58658 => x"082082",
   58659 => x"082082",
   58660 => x"082082",
   58661 => x"082082",
   58662 => x"082082",
   58663 => x"082082",
   58664 => x"082082",
   58665 => x"082082",
   58666 => x"082082",
   58667 => x"082082",
   58668 => x"082082",
   58669 => x"082082",
   58670 => x"082082",
   58671 => x"082082",
   58672 => x"082082",
   58673 => x"082082",
   58674 => x"082082",
   58675 => x"082082",
   58676 => x"082082",
   58677 => x"082082",
   58678 => x"082081",
   58679 => x"041041",
   58680 => x"041041",
   58681 => x"041041",
   58682 => x"041041",
   58683 => x"041041",
   58684 => x"041041",
   58685 => x"041041",
   58686 => x"041041",
   58687 => x"041041",
   58688 => x"041041",
   58689 => x"041041",
   58690 => x"041041",
   58691 => x"041041",
   58692 => x"041041",
   58693 => x"041041",
   58694 => x"041041",
   58695 => x"041041",
   58696 => x"041041",
   58697 => x"041041",
   58698 => x"041041",
   58699 => x"041041",
   58700 => x"041041",
   58701 => x"041041",
   58702 => x"041041",
   58703 => x"041000",
   58704 => x"000000",
   58705 => x"000000",
   58706 => x"000000",
   58707 => x"000000",
   58708 => x"000000",
   58709 => x"000abf",
   58710 => x"ffffff",
   58711 => x"ffffff",
   58712 => x"ffffff",
   58713 => x"ffffff",
   58714 => x"ffffff",
   58715 => x"ffffff",
   58716 => x"ffffff",
   58717 => x"ffffff",
   58718 => x"ffffff",
   58719 => x"ffffff",
   58720 => x"540000",
   58721 => x"000000",
   58722 => x"000000",
   58723 => x"000000",
   58724 => x"000000",
   58725 => x"000000",
   58726 => x"000000",
   58727 => x"000000",
   58728 => x"000000",
   58729 => x"000000",
   58730 => x"000000",
   58731 => x"000000",
   58732 => x"000000",
   58733 => x"000000",
   58734 => x"000000",
   58735 => x"000000",
   58736 => x"000000",
   58737 => x"000000",
   58738 => x"000000",
   58739 => x"000000",
   58740 => x"000000",
   58741 => x"000000",
   58742 => x"000000",
   58743 => x"000000",
   58744 => x"000000",
   58745 => x"000000",
   58746 => x"000000",
   58747 => x"000000",
   58748 => x"000000",
   58749 => x"000000",
   58750 => x"000000",
   58751 => x"000000",
   58752 => x"000000",
   58753 => x"000000",
   58754 => x"000000",
   58755 => x"000000",
   58756 => x"000000",
   58757 => x"000000",
   58758 => x"000000",
   58759 => x"000000",
   58760 => x"000000",
   58761 => x"000000",
   58762 => x"000000",
   58763 => x"000000",
   58764 => x"000000",
   58765 => x"000000",
   58766 => x"000000",
   58767 => x"000000",
   58768 => x"000000",
   58769 => x"000000",
   58770 => x"000000",
   58771 => x"000000",
   58772 => x"000000",
   58773 => x"000000",
   58774 => x"000000",
   58775 => x"000000",
   58776 => x"000000",
   58777 => x"000000",
   58778 => x"000000",
   58779 => x"000000",
   58780 => x"000000",
   58781 => x"000000",
   58782 => x"000000",
   58783 => x"000000",
   58784 => x"000000",
   58785 => x"000000",
   58786 => x"000000",
   58787 => x"000000",
   58788 => x"000000",
   58789 => x"000015",
   58790 => x"abffff",
   58791 => x"ffffff",
   58792 => x"ffffff",
   58793 => x"ffffff",
   58794 => x"ffffff",
   58795 => x"ffffff",
   58796 => x"ffffff",
   58797 => x"ffffff",
   58798 => x"ffffff",
   58799 => x"ffffff",
   58800 => x"ffffff",
   58801 => x"ffffff",
   58802 => x"ffffff",
   58803 => x"ffffff",
   58804 => x"ffffff",
   58805 => x"ffffff",
   58806 => x"ffffff",
   58807 => x"ffffff",
   58808 => x"ffffff",
   58809 => x"ffffff",
   58810 => x"ffffff",
   58811 => x"ffffff",
   58812 => x"ffffff",
   58813 => x"ffffff",
   58814 => x"ffffff",
   58815 => x"ffffff",
   58816 => x"ffffff",
   58817 => x"ffffff",
   58818 => x"ffffff",
   58819 => x"ffffff",
   58820 => x"ffffff",
   58821 => x"ffffff",
   58822 => x"ffffff",
   58823 => x"ffffff",
   58824 => x"ffffff",
   58825 => x"ffffff",
   58826 => x"ffffff",
   58827 => x"ffffff",
   58828 => x"ffffff",
   58829 => x"ffffff",
   58830 => x"ffffff",
   58831 => x"ffffff",
   58832 => x"ffffff",
   58833 => x"ffffff",
   58834 => x"ffffff",
   58835 => x"ffffff",
   58836 => x"ffffff",
   58837 => x"ffffff",
   58838 => x"ffffff",
   58839 => x"ffffff",
   58840 => x"ffffff",
   58841 => x"ffffff",
   58842 => x"ffffff",
   58843 => x"ffffff",
   58844 => x"ffffff",
   58845 => x"ffffff",
   58846 => x"ffffff",
   58847 => x"ffffff",
   58848 => x"ffffff",
   58849 => x"ffffff",
   58850 => x"ffffff",
   58851 => x"ffffff",
   58852 => x"ffffff",
   58853 => x"ffffff",
   58854 => x"ffffff",
   58855 => x"ffffff",
   58856 => x"ffffff",
   58857 => x"ffffff",
   58858 => x"ffffff",
   58859 => x"ffffff",
   58860 => x"ffffff",
   58861 => x"ffffff",
   58862 => x"ffffff",
   58863 => x"ffffff",
   58864 => x"ffffff",
   58865 => x"ffffff",
   58866 => x"ffffff",
   58867 => x"ffffff",
   58868 => x"ffffff",
   58869 => x"ffffff",
   58870 => x"ffffff",
   58871 => x"ffffff",
   58872 => x"ffffff",
   58873 => x"ffffff",
   58874 => x"ffffff",
   58875 => x"ffffff",
   58876 => x"ffffff",
   58877 => x"ffffff",
   58878 => x"ffffff",
   58879 => x"ffffff",
   58880 => x"ffffff",
   58881 => x"ffffff",
   58882 => x"ffffff",
   58883 => x"ffffff",
   58884 => x"ffffff",
   58885 => x"ffffff",
   58886 => x"ffffff",
   58887 => x"ffffff",
   58888 => x"ffffff",
   58889 => x"ffffff",
   58890 => x"ffffff",
   58891 => x"ffffff",
   58892 => x"ffffff",
   58893 => x"ffffff",
   58894 => x"ffffff",
   58895 => x"ffffff",
   58896 => x"ffffff",
   58897 => x"ffffff",
   58898 => x"ffffff",
   58899 => x"ffffff",
   58900 => x"ffffff",
   58901 => x"ffffff",
   58902 => x"ffffff",
   58903 => x"ffffff",
   58904 => x"ffffff",
   58905 => x"ffffff",
   58906 => x"ffffff",
   58907 => x"ffffff",
   58908 => x"ffffff",
   58909 => x"ffffff",
   58910 => x"ffffff",
   58911 => x"ffffff",
   58912 => x"ffffff",
   58913 => x"ffffff",
   58914 => x"ffffff",
   58915 => x"ffffff",
   58916 => x"ffffff",
   58917 => x"ffffff",
   58918 => x"ffffff",
   58919 => x"ffffff",
   58920 => x"ffffff",
   58921 => x"ffffff",
   58922 => x"ffffff",
   58923 => x"ffffff",
   58924 => x"ffffff",
   58925 => x"ffffff",
   58926 => x"ffffff",
   58927 => x"ffffff",
   58928 => x"ffffff",
   58929 => x"ffffff",
   58930 => x"ffffff",
   58931 => x"ffffff",
   58932 => x"ffffff",
   58933 => x"ffffff",
   58934 => x"ffffff",
   58935 => x"ffffff",
   58936 => x"ffffff",
   58937 => x"ffffff",
   58938 => x"ffffff",
   58939 => x"ffffff",
   58940 => x"ffffff",
   58941 => x"ffffff",
   58942 => x"ffffff",
   58943 => x"ffffff",
   58944 => x"ffffff",
   58945 => x"ffffff",
   58946 => x"ffffff",
   58947 => x"ffffff",
   58948 => x"ffffff",
   58949 => x"ffffff",
   58950 => x"ffffff",
   58951 => x"ffffff",
   58952 => x"ffffff",
   58953 => x"ffffff",
   58954 => x"ffffff",
   58955 => x"ffffff",
   58956 => x"ffffff",
   58957 => x"ffffff",
   58958 => x"ffffff",
   58959 => x"ffffff",
   58960 => x"ffffff",
   58961 => x"ffffff",
   58962 => x"ffffff",
   58963 => x"ffffff",
   58964 => x"ffffff",
   58965 => x"ffffff",
   58966 => x"ffffff",
   58967 => x"ffffff",
   58968 => x"ffffff",
   58969 => x"ffffff",
   58970 => x"ffffff",
   58971 => x"ffffff",
   58972 => x"ffffff",
   58973 => x"ffffff",
   58974 => x"ffffff",
   58975 => x"ffffff",
   58976 => x"ffffff",
   58977 => x"ffffff",
   58978 => x"ffffff",
   58979 => x"ffffff",
   58980 => x"ffffff",
   58981 => x"ffffff",
   58982 => x"ffffff",
   58983 => x"ffffff",
   58984 => x"ffffff",
   58985 => x"ffffff",
   58986 => x"ffffff",
   58987 => x"ffffff",
   58988 => x"ffffff",
   58989 => x"ffffff",
   58990 => x"ffffff",
   58991 => x"ffffff",
   58992 => x"ffffff",
   58993 => x"ffffff",
   58994 => x"ffffff",
   58995 => x"ffffff",
   58996 => x"ffffff",
   58997 => x"ffffff",
   58998 => x"ffffff",
   58999 => x"ffffff",
   59000 => x"ffffff",
   59001 => x"ffffff",
   59002 => x"ffffff",
   59003 => x"ffffff",
   59004 => x"ffffff",
   59005 => x"ffffff",
   59006 => x"ffffff",
   59007 => x"ffffff",
   59008 => x"ffffff",
   59009 => x"ffffff",
   59010 => x"ffffff",
   59011 => x"ffffff",
   59012 => x"ffffff",
   59013 => x"ffffff",
   59014 => x"ffffff",
   59015 => x"ffffff",
   59016 => x"ffffff",
   59017 => x"ffffff",
   59018 => x"ffffff",
   59019 => x"ffffff",
   59020 => x"ffffff",
   59021 => x"ffffff",
   59022 => x"ffffff",
   59023 => x"ffffff",
   59024 => x"ffffff",
   59025 => x"ffffff",
   59026 => x"ffffff",
   59027 => x"ffffff",
   59028 => x"ffffff",
   59029 => x"ffffff",
   59030 => x"ffffff",
   59031 => x"ffffff",
   59032 => x"ffffff",
   59033 => x"ffffff",
   59034 => x"ffffff",
   59035 => x"ffffff",
   59036 => x"ffffff",
   59037 => x"ffffff",
   59038 => x"ffffff",
   59039 => x"ffffff",
   59040 => x"ffffff",
   59041 => x"ffffff",
   59042 => x"ffffff",
   59043 => x"ffffff",
   59044 => x"ffffff",
   59045 => x"ffffff",
   59046 => x"ffffff",
   59047 => x"ffffff",
   59048 => x"ffffff",
   59049 => x"ffffff",
   59050 => x"ffffff",
   59051 => x"ffffff",
   59052 => x"ffffff",
   59053 => x"ffffff",
   59054 => x"ffffff",
   59055 => x"ffffff",
   59056 => x"ffffff",
   59057 => x"ffffff",
   59058 => x"ffffff",
   59059 => x"ffffff",
   59060 => x"ffffff",
   59061 => x"ffffff",
   59062 => x"ffffff",
   59063 => x"ffffff",
   59064 => x"ffffff",
   59065 => x"ffffff",
   59066 => x"ffffff",
   59067 => x"ffffff",
   59068 => x"ffffff",
   59069 => x"ffffff",
   59070 => x"ffffff",
   59071 => x"ffffff",
   59072 => x"ffffff",
   59073 => x"ffffff",
   59074 => x"ffffff",
   59075 => x"ffffff",
   59076 => x"ffffff",
   59077 => x"ffffff",
   59078 => x"ffffff",
   59079 => x"ffffff",
   59080 => x"ffffff",
   59081 => x"ffffff",
   59082 => x"ffffff",
   59083 => x"ffffff",
   59084 => x"ffffff",
   59085 => x"ffffff",
   59086 => x"ffffff",
   59087 => x"ffffff",
   59088 => x"ffffff",
   59089 => x"ffffff",
   59090 => x"ffffff",
   59091 => x"ffffff",
   59092 => x"ffffff",
   59093 => x"ffffff",
   59094 => x"ffffff",
   59095 => x"ffffff",
   59096 => x"ffffff",
   59097 => x"ffffff",
   59098 => x"ffffff",
   59099 => x"ffffff",
   59100 => x"ffffff",
   59101 => x"ffffff",
   59102 => x"ffffff",
   59103 => x"ffffff",
   59104 => x"ffffff",
   59105 => x"ffffff",
   59106 => x"ffffff",
   59107 => x"ffffff",
   59108 => x"ffffff",
   59109 => x"ffffff",
   59110 => x"ffffff",
   59111 => x"ffffff",
   59112 => x"ffffff",
   59113 => x"ffffff",
   59114 => x"ffffff",
   59115 => x"ffffff",
   59116 => x"ffffff",
   59117 => x"ffffff",
   59118 => x"ffffff",
   59119 => x"ffffff",
   59120 => x"ffffff",
   59121 => x"ffffff",
   59122 => x"ffffff",
   59123 => x"ffffff",
   59124 => x"ffffff",
   59125 => x"ffffff",
   59126 => x"ffffff",
   59127 => x"ffffff",
   59128 => x"ffffff",
   59129 => x"ffffff",
   59130 => x"ffffff",
   59131 => x"ffffff",
   59132 => x"ffffff",
   59133 => x"ffffff",
   59134 => x"ffffff",
   59135 => x"ffffff",
   59136 => x"ffffff",
   59137 => x"ffffff",
   59138 => x"ffffff",
   59139 => x"ffffff",
   59140 => x"ffffff",
   59141 => x"ffffff",
   59142 => x"ffffff",
   59143 => x"ffffff",
   59144 => x"ffffff",
   59145 => x"ffffff",
   59146 => x"ffffff",
   59147 => x"ffffff",
   59148 => x"ffffff",
   59149 => x"ffffff",
   59150 => x"ffffff",
   59151 => x"ffffff",
   59152 => x"ffffff",
   59153 => x"ffffff",
   59154 => x"ffffff",
   59155 => x"ffffff",
   59156 => x"ffffff",
   59157 => x"ffffff",
   59158 => x"ffffff",
   59159 => x"ffffff",
   59160 => x"ffffff",
   59161 => x"ffffff",
   59162 => x"ffffff",
   59163 => x"ffffff",
   59164 => x"ffffff",
   59165 => x"ffffff",
   59166 => x"ffffff",
   59167 => x"ffffff",
   59168 => x"ffffff",
   59169 => x"ffffff",
   59170 => x"ffffff",
   59171 => x"ffffff",
   59172 => x"ffffff",
   59173 => x"ffffff",
   59174 => x"ffffff",
   59175 => x"ffffff",
   59176 => x"ffffff",
   59177 => x"ffffff",
   59178 => x"ffffff",
   59179 => x"ffffff",
   59180 => x"ffffff",
   59181 => x"ffffff",
   59182 => x"ffffff",
   59183 => x"ffffff",
   59184 => x"ffffff",
   59185 => x"ffffff",
   59186 => x"ffffff",
   59187 => x"ffffff",
   59188 => x"ffffff",
   59189 => x"ffffff",
   59190 => x"ffffff",
   59191 => x"ffffff",
   59192 => x"ffffff",
   59193 => x"ffffff",
   59194 => x"ffffff",
   59195 => x"ffffff",
   59196 => x"ffffff",
   59197 => x"ffffff",
   59198 => x"ffffff",
   59199 => x"ffffff",
   59200 => x"ffffff",
   59201 => x"ffffff",
   59202 => x"ffffff",
   59203 => x"ffffff",
   59204 => x"ffffff",
   59205 => x"ffffff",
   59206 => x"ffffff",
   59207 => x"ffffff",
   59208 => x"ffffff",
   59209 => x"ffffff",
   59210 => x"ffffff",
   59211 => x"ffffff",
   59212 => x"ffffff",
   59213 => x"ffffff",
   59214 => x"ffffff",
   59215 => x"ffffff",
   59216 => x"ffffff",
   59217 => x"ffffff",
   59218 => x"ffffff",
   59219 => x"ffffff",
   59220 => x"ffffff",
   59221 => x"ffffff",
   59222 => x"ffffff",
   59223 => x"ffffff",
   59224 => x"ffffff",
   59225 => x"ffffff",
   59226 => x"ffffff",
   59227 => x"ffffff",
   59228 => x"ffffff",
   59229 => x"ffffff",
   59230 => x"ffffff",
   59231 => x"ffffff",
   59232 => x"ffffff",
   59233 => x"ffffff",
   59234 => x"ffffff",
   59235 => x"ffffff",
   59236 => x"ffffff",
   59237 => x"ffffff",
   59238 => x"ffffff",
   59239 => x"ffffff",
   59240 => x"ffffff",
   59241 => x"ffffff",
   59242 => x"ffffff",
   59243 => x"ffffff",
   59244 => x"ffffff",
   59245 => x"ffffff",
   59246 => x"ffffff",
   59247 => x"ffffff",
   59248 => x"ffffff",
   59249 => x"ffffff",
   59250 => x"ffffff",
   59251 => x"ffffff",
   59252 => x"ffffff",
   59253 => x"ffffff",
   59254 => x"ffffff",
   59255 => x"ffffff",
   59256 => x"ffffff",
   59257 => x"ffffff",
   59258 => x"ffffff",
   59259 => x"ffffff",
   59260 => x"ffffff",
   59261 => x"ffffff",
   59262 => x"ffffff",
   59263 => x"ffffff",
   59264 => x"ffffff",
   59265 => x"ffffff",
   59266 => x"ffffff",
   59267 => x"ffffff",
   59268 => x"ffffff",
   59269 => x"ffffff",
   59270 => x"ffffff",
   59271 => x"ffffff",
   59272 => x"ffffff",
   59273 => x"ffffff",
   59274 => x"ffffff",
   59275 => x"ffffff",
   59276 => x"ffffff",
   59277 => x"ffffff",
   59278 => x"ffffff",
   59279 => x"ffffff",
   59280 => x"ffffff",
   59281 => x"ffffff",
   59282 => x"ffffff",
   59283 => x"ffffff",
   59284 => x"ffffff",
   59285 => x"ffffff",
   59286 => x"ffffff",
   59287 => x"ffffff",
   59288 => x"ffffff",
   59289 => x"ffffff",
   59290 => x"ffffff",
   59291 => x"ffffff",
   59292 => x"ffffff",
   59293 => x"ffffff",
   59294 => x"ffffff",
   59295 => x"ffffff",
   59296 => x"ffffff",
   59297 => x"ffffff",
   59298 => x"ffffff",
   59299 => x"ffffff",
   59300 => x"ffffff",
   59301 => x"ffffff",
   59302 => x"ffffff",
   59303 => x"ffffff",
   59304 => x"ffffff",
   59305 => x"ffffff",
   59306 => x"ffffff",
   59307 => x"ffffff",
   59308 => x"ffffff",
   59309 => x"ffffff",
   59310 => x"ffffff",
   59311 => x"ffffff",
   59312 => x"ffffff",
   59313 => x"ffffff",
   59314 => x"ffffff",
   59315 => x"ffffff",
   59316 => x"ffffff",
   59317 => x"ffffff",
   59318 => x"ffffff",
   59319 => x"ffffff",
   59320 => x"ffffff",
   59321 => x"ffffff",
   59322 => x"ffffff",
   59323 => x"ffffff",
   59324 => x"ffffff",
   59325 => x"ffffff",
   59326 => x"ffffff",
   59327 => x"ffffff",
   59328 => x"ffffff",
   59329 => x"ffffff",
   59330 => x"ffffff",
   59331 => x"ffffff",
   59332 => x"ffffff",
   59333 => x"ffffff",
   59334 => x"ffffff",
   59335 => x"ffffff",
   59336 => x"ffffff",
   59337 => x"ffffff",
   59338 => x"ffffff",
   59339 => x"ffffff",
   59340 => x"ffffff",
   59341 => x"ffffff",
   59342 => x"ffffff",
   59343 => x"ffffff",
   59344 => x"ffffff",
   59345 => x"ffffff",
   59346 => x"ffffff",
   59347 => x"ffffff",
   59348 => x"ffffff",
   59349 => x"ffffff",
   59350 => x"ffffff",
   59351 => x"ffffff",
   59352 => x"ffffff",
   59353 => x"ffffff",
   59354 => x"ffffff",
   59355 => x"ffffff",
   59356 => x"ffffff",
   59357 => x"ffffff",
   59358 => x"ffffff",
   59359 => x"ffffff",
   59360 => x"ffffff",
   59361 => x"ffffff",
   59362 => x"ffffff",
   59363 => x"ffffff",
   59364 => x"ffffff",
   59365 => x"ffffff",
   59366 => x"ffffff",
   59367 => x"ffffff",
   59368 => x"ffffff",
   59369 => x"ffffff",
   59370 => x"ffffff",
   59371 => x"ffffff",
   59372 => x"ffffff",
   59373 => x"ffffff",
   59374 => x"ffffff",
   59375 => x"ffffff",
   59376 => x"ffffff",
   59377 => x"ffffff",
   59378 => x"ffffff",
   59379 => x"ffffff",
   59380 => x"ffffff",
   59381 => x"ffffff",
   59382 => x"ffffff",
   59383 => x"ffffff",
   59384 => x"ffffff",
   59385 => x"ffffff",
   59386 => x"ffffff",
   59387 => x"ffffff",
   59388 => x"ffffff",
   59389 => x"ffffff",
   59390 => x"ffffff",
   59391 => x"ffffff",
   59392 => x"ffffff",
   59393 => x"ffffff",
   59394 => x"ffffff",
   59395 => x"ffffff",
   59396 => x"ffffff",
   59397 => x"ffffff",
   59398 => x"ffffff",
   59399 => x"ffffff",
   59400 => x"ffffff",
   59401 => x"ffffff",
   59402 => x"ffffff",
   59403 => x"ffffff",
   59404 => x"ffffff",
   59405 => x"ffffff",
   59406 => x"ffffff",
   59407 => x"ffffff",
   59408 => x"ffffff",
   59409 => x"ffffff",
   59410 => x"ffffff",
   59411 => x"ffffff",
   59412 => x"ffffff",
   59413 => x"ffffff",
   59414 => x"ffffff",
   59415 => x"ffffff",
   59416 => x"ffffff",
   59417 => x"ffffff",
   59418 => x"ffffff",
   59419 => x"ffffff",
   59420 => x"ffffff",
   59421 => x"ffffff",
   59422 => x"ffffff",
   59423 => x"ffffff",
   59424 => x"ffffff",
   59425 => x"ffffff",
   59426 => x"ffffff",
   59427 => x"ffffff",
   59428 => x"ffffff",
   59429 => x"ffffff",
   59430 => x"ffffff",
   59431 => x"ffffff",
   59432 => x"ffffff",
   59433 => x"ffffff",
   59434 => x"ffffff",
   59435 => x"ffffff",
   59436 => x"ffffff",
   59437 => x"ffffff",
   59438 => x"ffffff",
   59439 => x"ffffff",
   59440 => x"ffffff",
   59441 => x"ffffff",
   59442 => x"ffffff",
   59443 => x"ffffff",
   59444 => x"ffffff",
   59445 => x"ffffff",
   59446 => x"ffffff",
   59447 => x"ffffff",
   59448 => x"ffffff",
   59449 => x"ffffff",
   59450 => x"ffffff",
   59451 => x"ffffff",
   59452 => x"ffffff",
   59453 => x"ffffff",
   59454 => x"ffffff",
   59455 => x"ffffff",
   59456 => x"ffffff",
   59457 => x"ffffff",
   59458 => x"ffffff",
   59459 => x"ffffff",
   59460 => x"ffffff",
   59461 => x"ffffff",
   59462 => x"ffffff",
   59463 => x"ffffff",
   59464 => x"ffffff",
   59465 => x"ffffff",
   59466 => x"ffffff",
   59467 => x"ffffff",
   59468 => x"ffffff",
   59469 => x"ffffff",
   59470 => x"ffffff",
   59471 => x"ffffff",
   59472 => x"ffffff",
   59473 => x"ffffff",
   59474 => x"ffffff",
   59475 => x"ffffff",
   59476 => x"ffffff",
   59477 => x"ffffff",
   59478 => x"ffffff",
   59479 => x"ffffff",
   59480 => x"ffffff",
   59481 => x"ffffff",
   59482 => x"ffffff",
   59483 => x"ffffff",
   59484 => x"ffffff",
   59485 => x"ffffff",
   59486 => x"ffffff",
   59487 => x"ffffff",
   59488 => x"ffffff",
   59489 => x"ffffff",
   59490 => x"ffffff",
   59491 => x"ffffff",
   59492 => x"ffffff",
   59493 => x"ffffff",
   59494 => x"ffffff",
   59495 => x"ffffff",
   59496 => x"ffffff",
   59497 => x"ffffff",
   59498 => x"ffffff",
   59499 => x"ffffff",
   59500 => x"ffffff",
   59501 => x"ffffff",
   59502 => x"ffffff",
   59503 => x"ffffff",
   59504 => x"ffffff",
   59505 => x"ffffff",
   59506 => x"ffffff",
   59507 => x"ffffff",
   59508 => x"ffffff",
   59509 => x"ffffff",
   59510 => x"ffffff",
   59511 => x"ffffff",
   59512 => x"ffffff",
   59513 => x"ffffff",
   59514 => x"ffffff",
   59515 => x"ffffff",
   59516 => x"ffffff",
   59517 => x"ffffff",
   59518 => x"ffffff",
   59519 => x"ffffff",
   59520 => x"ffffff",
   59521 => x"ffffff",
   59522 => x"ffffff",
   59523 => x"ffffff",
   59524 => x"ffffff",
   59525 => x"ffffff",
   59526 => x"ffffff",
   59527 => x"ffffff",
   59528 => x"ffffff",
   59529 => x"ffffff",
   59530 => x"ffffff",
   59531 => x"ffffff",
   59532 => x"ffffff",
   59533 => x"ffffff",
   59534 => x"ffffff",
   59535 => x"ffffff",
   59536 => x"ffffff",
   59537 => x"ffffff",
   59538 => x"ffffff",
   59539 => x"ffffff",
   59540 => x"ffffff",
   59541 => x"ffffff",
   59542 => x"ffffff",
   59543 => x"ffffff",
   59544 => x"ffffff",
   59545 => x"ffffff",
   59546 => x"ffffff",
   59547 => x"ffffff",
   59548 => x"ffffff",
   59549 => x"ffffff",
   59550 => x"ffffff",
   59551 => x"ffffff",
   59552 => x"ffffff",
   59553 => x"ffffff",
   59554 => x"ffffff",
   59555 => x"ffffff",
   59556 => x"ffffff",
   59557 => x"ffffff",
   59558 => x"ffffff",
   59559 => x"ffffff",
   59560 => x"ffffff",
   59561 => x"ffffff",
   59562 => x"ffffff",
   59563 => x"ffffff",
   59564 => x"ffffff",
   59565 => x"ffffff",
   59566 => x"ffffff",
   59567 => x"ffffff",
   59568 => x"ffffff",
   59569 => x"ffffff",
   59570 => x"ffffff",
   59571 => x"ffffff",
   59572 => x"ffffff",
   59573 => x"ffffff",
   59574 => x"ffffff",
   59575 => x"ffffff",
   59576 => x"ffffff",
   59577 => x"ffffff",
   59578 => x"ffffff",
   59579 => x"ffffff",
   59580 => x"ffffff",
   59581 => x"ffffff",
   59582 => x"ffffff",
   59583 => x"ffffff",
   59584 => x"ffffff",
   59585 => x"ffffff",
   59586 => x"ffffff",
   59587 => x"ffffff",
   59588 => x"ffffff",
   59589 => x"ffffff",
   59590 => x"ffffff",
   59591 => x"ffffff",
   59592 => x"ffffff",
   59593 => x"ffffff",
   59594 => x"ffffff",
   59595 => x"ffffff",
   59596 => x"ffffff",
   59597 => x"ffffff",
   59598 => x"ffffff",
   59599 => x"ffffff",
   59600 => x"ffffff",
   59601 => x"ffffff",
   59602 => x"ffffff",
   59603 => x"ffffff",
   59604 => x"ffffff",
   59605 => x"ffffff",
   59606 => x"ffffff",
   59607 => x"ffffff",
   59608 => x"ffffff",
   59609 => x"ffffff",
   59610 => x"ffffff",
   59611 => x"ffffff",
   59612 => x"ffffff",
   59613 => x"ffffff",
   59614 => x"ffffff",
   59615 => x"ffffff",
   59616 => x"ffffff",
   59617 => x"ffffff",
   59618 => x"ffffff",
   59619 => x"ffffff",
   59620 => x"ffffff",
   59621 => x"ffffff",
   59622 => x"ffffff",
   59623 => x"ffffff",
   59624 => x"ffffff",
   59625 => x"ffffff",
   59626 => x"ffffff",
   59627 => x"ffffff",
   59628 => x"ffffff",
   59629 => x"ffffff",
   59630 => x"ffffff",
   59631 => x"ffffff",
   59632 => x"ffffff",
   59633 => x"ffffff",
   59634 => x"ffffff",
   59635 => x"ffffff",
   59636 => x"ffffff",
   59637 => x"ffffff",
   59638 => x"ffffff",
   59639 => x"ffffff",
   59640 => x"ffffff",
   59641 => x"ffffff",
   59642 => x"ffffff",
   59643 => x"ffffff",
   59644 => x"ffffff",
   59645 => x"ffffff",
   59646 => x"ffffff",
   59647 => x"ffffff",
   59648 => x"ffffff",
   59649 => x"ffffff",
   59650 => x"ffffff",
   59651 => x"ffffff",
   59652 => x"ffffff",
   59653 => x"ffffff",
   59654 => x"ffffff",
   59655 => x"ffffff",
   59656 => x"ffffff",
   59657 => x"ffffff",
   59658 => x"ffffff",
   59659 => x"ffffff",
   59660 => x"ffffff",
   59661 => x"ffffff",
   59662 => x"ffffff",
   59663 => x"ffffff",
   59664 => x"ffffff",
   59665 => x"ffffff",
   59666 => x"ffffff",
   59667 => x"ffffff",
   59668 => x"ffffff",
   59669 => x"ffffff",
   59670 => x"ffffff",
   59671 => x"ffffff",
   59672 => x"ffffff",
   59673 => x"ffffff",
   59674 => x"ffffff",
   59675 => x"ffffff",
   59676 => x"ffffff",
   59677 => x"ffffff",
   59678 => x"ffffff",
   59679 => x"ffffff",
   59680 => x"ffffff",
   59681 => x"ffffff",
   59682 => x"ffffff",
   59683 => x"ffffff",
   59684 => x"ffffff",
   59685 => x"ffffff",
   59686 => x"ffffff",
   59687 => x"ffffff",
   59688 => x"ffffff",
   59689 => x"ffffff",
   59690 => x"ffffff",
   59691 => x"ffffff",
   59692 => x"ffffff",
   59693 => x"ffffff",
   59694 => x"ffffff",
   59695 => x"ffffff",
   59696 => x"ffffff",
   59697 => x"ffffff",
   59698 => x"ffffff",
   59699 => x"ffffff",
   59700 => x"ffffff",
   59701 => x"ffffff",
   59702 => x"ffffff",
   59703 => x"ffffff",
   59704 => x"ffffff",
   59705 => x"ffffff",
   59706 => x"ffffff",
   59707 => x"ffffff",
   59708 => x"ffffff",
   59709 => x"ffffff",
   59710 => x"ffffff",
   59711 => x"ffffff",
   59712 => x"ffffff",
   59713 => x"ffffff",
   59714 => x"ffffff",
   59715 => x"ffffff",
   59716 => x"ffffff",
   59717 => x"ffffff",
   59718 => x"ffffff",
   59719 => x"ffffff",
   59720 => x"ffffff",
   59721 => x"ffffff",
   59722 => x"ffffff",
   59723 => x"ffffff",
   59724 => x"ffffff",
   59725 => x"ffffff",
   59726 => x"ffffff",
   59727 => x"ffffff",
   59728 => x"ffffff",
   59729 => x"ffffff",
   59730 => x"ffffff",
   59731 => x"ffffff",
   59732 => x"ffffff",
   59733 => x"ffffff",
   59734 => x"ffffff",
   59735 => x"ffffff",
   59736 => x"ffffff",
   59737 => x"ffffff",
   59738 => x"ffffff",
   59739 => x"ffffff",
   59740 => x"ffffff",
   59741 => x"ffffff",
   59742 => x"ffffff",
   59743 => x"ffffff",
   59744 => x"ffffff",
   59745 => x"ffffff",
   59746 => x"ffffff",
   59747 => x"ffffff",
   59748 => x"ffffff",
   59749 => x"ffffff",
   59750 => x"ffffff",
   59751 => x"ffffff",
   59752 => x"ffffff",
   59753 => x"ffffff",
   59754 => x"ffffff",
   59755 => x"ffffff",
   59756 => x"ffffff",
   59757 => x"ffffff",
   59758 => x"ffffff",
   59759 => x"ffffff",
   59760 => x"ffffff",
   59761 => x"ffffff",
   59762 => x"ffffff",
   59763 => x"ffffff",
   59764 => x"ffffff",
   59765 => x"ffffff",
   59766 => x"ffffff",
   59767 => x"ffffff",
   59768 => x"ffffff",
   59769 => x"ffffff",
   59770 => x"ffffff",
   59771 => x"ffffff",
   59772 => x"ffffff",
   59773 => x"ffffff",
   59774 => x"ffffff",
   59775 => x"ffffff",
   59776 => x"ffffff",
   59777 => x"ffffff",
   59778 => x"ffffff",
   59779 => x"ffffff",
   59780 => x"ffffff",
   59781 => x"ffffff",
   59782 => x"ffffff",
   59783 => x"ffffff",
   59784 => x"ffffff",
   59785 => x"ffffff",
   59786 => x"ffffff",
   59787 => x"ffffff",
   59788 => x"ffffff",
   59789 => x"ffffff",
   59790 => x"ffffff",
   59791 => x"ffffff",
   59792 => x"ffffff",
   59793 => x"ffffff",
   59794 => x"ffffff",
   59795 => x"ffffff",
   59796 => x"ffffff",
   59797 => x"ffffff",
   59798 => x"ffffff",
   59799 => x"ffffff",
   59800 => x"ffffff",
   59801 => x"ffffff",
   59802 => x"ffffff",
   59803 => x"ffffff",
   59804 => x"ffffff",
   59805 => x"ffffff",
   59806 => x"ffffff",
   59807 => x"ffffff",
   59808 => x"ffffff",
   59809 => x"ffffff",
   59810 => x"ffffff",
   59811 => x"ffffff",
   59812 => x"ffffff",
   59813 => x"ffffff",
   59814 => x"ffffff",
   59815 => x"ffffff",
   59816 => x"ffffff",
   59817 => x"ffffff",
   59818 => x"ffffff",
   59819 => x"ffffff",
   59820 => x"ffffff",
   59821 => x"ffffff",
   59822 => x"ffffff",
   59823 => x"ffffff",
   59824 => x"ffffff",
   59825 => x"ffffff",
   59826 => x"ffffff",
   59827 => x"ffffff",
   59828 => x"ffffff",
   59829 => x"ffffff",
   59830 => x"ffffff",
   59831 => x"ffffff",
   59832 => x"ffffff",
   59833 => x"ffffff",
   59834 => x"ffffff",
   59835 => x"ffffff",
   59836 => x"ffffff",
   59837 => x"ffffff",
   59838 => x"ffffff",
   59839 => x"ffffff",
   59840 => x"ffffff",
   59841 => x"ffffff",
   59842 => x"ffffff",
   59843 => x"ffffff",
   59844 => x"ffffff",
   59845 => x"ffffff",
   59846 => x"ffffff",
   59847 => x"ffffff",
   59848 => x"ffffff",
   59849 => x"ffffff",
   59850 => x"ffffff",
   59851 => x"ffffff",
   59852 => x"ffffff",
   59853 => x"ffffff",
   59854 => x"ffffff",
   59855 => x"ffffff",
   59856 => x"ffffff",
   59857 => x"ffffff",
   59858 => x"ffffff",
   59859 => x"ffffff",
   59860 => x"ffffff",
   59861 => x"ffffff",
   59862 => x"ffffff",
   59863 => x"ffffff",
   59864 => x"ffffff",
   59865 => x"ffffff",
   59866 => x"ffffff",
   59867 => x"ffffff",
   59868 => x"ffffff",
   59869 => x"ffffff",
   59870 => x"ffffff",
   59871 => x"ffffff",
   59872 => x"ffffff",
   59873 => x"ffffff",
   59874 => x"ffffff",
   59875 => x"ffffff",
   59876 => x"ffffff",
   59877 => x"ffffff",
   59878 => x"ffffff",
   59879 => x"ffffff",
   59880 => x"ffffff",
   59881 => x"ffffff",
   59882 => x"ffffff",
   59883 => x"ffffff",
   59884 => x"ffffff",
   59885 => x"ffffff",
   59886 => x"ffffff",
   59887 => x"ffffff",
   59888 => x"ffffff",
   59889 => x"ffffff",
   59890 => x"ffffff",
   59891 => x"ffffff",
   59892 => x"ffffff",
   59893 => x"ffffff",
   59894 => x"ffffff",
   59895 => x"ffffff",
   59896 => x"ffffff",
   59897 => x"ffffff",
   59898 => x"ffffff",
   59899 => x"ffffff",
   59900 => x"ffffff",
   59901 => x"ffffff",
   59902 => x"ffffff",
   59903 => x"ffffff",
   59904 => x"ffffff",
   59905 => x"ffffff",
   59906 => x"ffffff",
   59907 => x"ffffff",
   59908 => x"ffffff",
   59909 => x"ffffff",
   59910 => x"ffffff",
   59911 => x"ffffff",
   59912 => x"ffffff",
   59913 => x"ffffff",
   59914 => x"ffffff",
   59915 => x"ffffff",
   59916 => x"ffffff",
   59917 => x"ffffff",
   59918 => x"ffffff",
   59919 => x"ffffff",
   59920 => x"ffffff",
   59921 => x"ffffff",
   59922 => x"ffffff",
   59923 => x"ffffff",
   59924 => x"ffffff",
   59925 => x"ffffff",
   59926 => x"ffffff",
   59927 => x"ffffff",
   59928 => x"ffffff",
   59929 => x"ffffff",
   59930 => x"ffffff",
   59931 => x"ffffff",
   59932 => x"ffffff",
   59933 => x"ffffff",
   59934 => x"ffffff",
   59935 => x"ffffff",
   59936 => x"ffffff",
   59937 => x"ffffff",
   59938 => x"ffffff",
   59939 => x"ffffff",
   59940 => x"ffffff",
   59941 => x"ffffff",
   59942 => x"ffffff",
   59943 => x"ffffff",
   59944 => x"ffffff",
   59945 => x"ffffff",
   59946 => x"ffffff",
   59947 => x"ffffff",
   59948 => x"ffffff",
   59949 => x"ffffff",
   59950 => x"ffffff",
   59951 => x"ffffff",
   59952 => x"ffffff",
   59953 => x"ffffff",
   59954 => x"ffffff",
   59955 => x"ffffff",
   59956 => x"ffffff",
   59957 => x"ffffff",
   59958 => x"ffffff",
   59959 => x"ffffff",
   59960 => x"ffffff",
   59961 => x"ffffff",
   59962 => x"ffffff",
   59963 => x"ffffff",
   59964 => x"ffffff",
   59965 => x"ffffff",
   59966 => x"ffffff",
   59967 => x"ffffff",
   59968 => x"ffffff",
   59969 => x"ffffff",
   59970 => x"ffffff",
   59971 => x"ffffff",
   59972 => x"ffffff",
   59973 => x"ffffff",
   59974 => x"ffffff",
   59975 => x"ffffff",
   59976 => x"ffffff",
   59977 => x"ffffff",
   59978 => x"ffffff",
   59979 => x"ffffff",
   59980 => x"ffffff",
   59981 => x"ffffff",
   59982 => x"ffffff",
   59983 => x"ffffff",
   59984 => x"ffffff",
   59985 => x"ffffff",
   59986 => x"ffffff",
   59987 => x"ffffff",
   59988 => x"ffffff",
   59989 => x"ffffff",
   59990 => x"ffffff",
   59991 => x"ffffff",
   59992 => x"ffffff",
   59993 => x"ffffff",
   59994 => x"ffffff",
   59995 => x"ffffff",
   59996 => x"ffffff",
   59997 => x"ffffff",
   59998 => x"ffffff",
   59999 => x"ffffff",
   60000 => x"ffffff",
   60001 => x"ffffff",
   60002 => x"ffffff",
   60003 => x"ffffff",
   60004 => x"ffffff",
   60005 => x"ffffff",
   60006 => x"ffffff",
   60007 => x"ffffff",
   60008 => x"ffffff",
   60009 => x"ffffff",
   60010 => x"ffffff",
   60011 => x"ffffff",
   60012 => x"ffffff",
   60013 => x"ffffff",
   60014 => x"ffffff",
   60015 => x"ffffff",
   60016 => x"ffffff",
   60017 => x"ffffff",
   60018 => x"ffffff",
   60019 => x"ffffff",
   60020 => x"ffffff",
   60021 => x"ffffff",
   60022 => x"ffffff",
   60023 => x"ffffff",
   60024 => x"ffffff",
   60025 => x"ffffff",
   60026 => x"ffffff",
   60027 => x"ffffff",
   60028 => x"ffffff",
   60029 => x"ffffff",
   60030 => x"ffffff",
   60031 => x"ffffff",
   60032 => x"ffffff",
   60033 => x"ffffff",
   60034 => x"ffffff",
   60035 => x"ffffff",
   60036 => x"ffffff",
   60037 => x"ffffff",
   60038 => x"ffffff",
   60039 => x"ffffff",
   60040 => x"ffffff",
   60041 => x"ffffff",
   60042 => x"ffffff",
   60043 => x"ffffff",
   60044 => x"ffffff",
   60045 => x"ffffff",
   60046 => x"ffffff",
   60047 => x"ffffff",
   60048 => x"ffffff",
   60049 => x"ffffff",
   60050 => x"ffffff",
   60051 => x"ffffff",
   60052 => x"ffffff",
   60053 => x"ffffff",
   60054 => x"ffffff",
   60055 => x"ffffff",
   60056 => x"ffffff",
   60057 => x"ffffff",
   60058 => x"ffffff",
   60059 => x"ffffff",
   60060 => x"ffffff",
   60061 => x"ffffff",
   60062 => x"ffffff",
   60063 => x"ffffff",
   60064 => x"ffffff",
   60065 => x"ffffff",
   60066 => x"ffffff",
   60067 => x"ffffff",
   60068 => x"ffffff",
   60069 => x"ffffff",
   60070 => x"ffffff",
   60071 => x"ffffff",
   60072 => x"ffffff",
   60073 => x"ffffff",
   60074 => x"ffffff",
   60075 => x"ffffff",
   60076 => x"ffffff",
   60077 => x"ffffff",
   60078 => x"ffffff",
   60079 => x"ffffff",
   60080 => x"ffffff",
   60081 => x"ffffff",
   60082 => x"ffffff",
   60083 => x"ffffff",
   60084 => x"ffffff",
   60085 => x"ffffff",
   60086 => x"ffffff",
   60087 => x"ffffff",
   60088 => x"ffffff",
   60089 => x"ffffff",
   60090 => x"ffffff",
   60091 => x"ffffff",
   60092 => x"ffffff",
   60093 => x"ffffff",
   60094 => x"ffffff",
   60095 => x"ffffff",
   60096 => x"ffffff",
   60097 => x"ffffff",
   60098 => x"ffffff",
   60099 => x"ffffff",
   60100 => x"ffffff",
   60101 => x"ffffff",
   60102 => x"ffffff",
   60103 => x"ffffff",
   60104 => x"ffffff",
   60105 => x"ffffff",
   60106 => x"ffffff",
   60107 => x"ffffff",
   60108 => x"ffffff",
   60109 => x"ffffff",
   60110 => x"ffffff",
   60111 => x"ffffff",
   60112 => x"ffffff",
   60113 => x"ffffff",
   60114 => x"ffffff",
   60115 => x"ffffff",
   60116 => x"ffffff",
   60117 => x"ffffff",
   60118 => x"ffffff",
   60119 => x"ffffff",
   60120 => x"ffffff",
   60121 => x"ffffff",
   60122 => x"ffffff",
   60123 => x"ffffff",
   60124 => x"ffffff",
   60125 => x"ffffff",
   60126 => x"ffffff",
   60127 => x"ffffff",
   60128 => x"ffffff",
   60129 => x"ffffff",
   60130 => x"ffffff",
   60131 => x"ffffff",
   60132 => x"ffffff",
   60133 => x"ffffff",
   60134 => x"ffffff",
   60135 => x"ffffff",
   60136 => x"ffffff",
   60137 => x"ffffff",
   60138 => x"ffffff",
   60139 => x"ffffff",
   60140 => x"ffffff",
   60141 => x"ffffff",
   60142 => x"ffffff",
   60143 => x"ffffff",
   60144 => x"ffffff",
   60145 => x"ffffff",
   60146 => x"ffffff",
   60147 => x"ffffff",
   60148 => x"ffffff",
   60149 => x"ffffff",
   60150 => x"ffffff",
   60151 => x"ffffff",
   60152 => x"ffffff",
   60153 => x"ffffff",
   60154 => x"ffffff",
   60155 => x"ffffff",
   60156 => x"ffffff",
   60157 => x"ffffff",
   60158 => x"ffffff",
   60159 => x"ffffff",
   60160 => x"ffffff",
   60161 => x"ffffff",
   60162 => x"ffffff",
   60163 => x"ffffff",
   60164 => x"ffffff",
   60165 => x"ffffff",
   60166 => x"ffffff",
   60167 => x"ffffff",
   60168 => x"ffffff",
   60169 => x"ffffff",
   60170 => x"ffffff",
   60171 => x"ffffff",
   60172 => x"ffffff",
   60173 => x"ffffff",
   60174 => x"ffffff",
   60175 => x"ffffff",
   60176 => x"ffffff",
   60177 => x"ffffff",
   60178 => x"ffffff",
   60179 => x"ffffff",
   60180 => x"ffffff",
   60181 => x"ffffff",
   60182 => x"ffffff",
   60183 => x"ffffff",
   60184 => x"ffffff",
   60185 => x"ffffff",
   60186 => x"ffffff",
   60187 => x"ffffff",
   60188 => x"ffffff",
   60189 => x"ffffff",
   60190 => x"ffffff",
   60191 => x"ffffff",
   60192 => x"ffffff",
   60193 => x"ffffff",
   60194 => x"ffffff",
   60195 => x"ffffff",
   60196 => x"ffffff",
   60197 => x"ffffff",
   60198 => x"ffffff",
   60199 => x"ffffff",
   60200 => x"ffffff",
   60201 => x"ffffff",
   60202 => x"ffffff",
   60203 => x"ffffff",
   60204 => x"ffffff",
   60205 => x"ffffff",
   60206 => x"ffffff",
   60207 => x"ffffff",
   60208 => x"ffffff",
   60209 => x"ffffff",
   60210 => x"ffffff",
   60211 => x"ffffff",
   60212 => x"ffffff",
   60213 => x"ffffff",
   60214 => x"ffffff",
   60215 => x"ffffff",
   60216 => x"ffffff",
   60217 => x"ffffff",
   60218 => x"ffffff",
   60219 => x"ffffff",
   60220 => x"ffffff",
   60221 => x"ffffff",
   60222 => x"ffffff",
   60223 => x"ffffff",
   60224 => x"ffffff",
   60225 => x"ffffff",
   60226 => x"ffffff",
   60227 => x"ffffff",
   60228 => x"ffffff",
   60229 => x"ffffff",
   60230 => x"ffffff",
   60231 => x"ffffff",
   60232 => x"ffffff",
   60233 => x"ffffff",
   60234 => x"ffffff",
   60235 => x"ffffff",
   60236 => x"ffffff",
   60237 => x"ffffff",
   60238 => x"ffffff",
   60239 => x"ffffff",
   60240 => x"ffffff",
   60241 => x"ffffff",
   60242 => x"ffffff",
   60243 => x"ffffff",
   60244 => x"ffffff",
   60245 => x"ffffff",
   60246 => x"ffffff",
   60247 => x"ffffff",
   60248 => x"ffffff",
   60249 => x"ffffff",
   60250 => x"ffffff",
   60251 => x"ffffff",
   60252 => x"ffffff",
   60253 => x"ffffff",
   60254 => x"ffffff",
   60255 => x"ffffff",
   60256 => x"ffffff",
   60257 => x"ffffff",
   60258 => x"ffffff",
   60259 => x"ffffff",
   60260 => x"ffffff",
   60261 => x"ffffff",
   60262 => x"ffffff",
   60263 => x"ffffff",
   60264 => x"ffffff",
   60265 => x"ffffff",
   60266 => x"ffffff",
   60267 => x"ffffff",
   60268 => x"ffffff",
   60269 => x"ffffff",
   60270 => x"ffffff",
   60271 => x"ffffff",
   60272 => x"ffffff",
   60273 => x"ffffff",
   60274 => x"ffffff",
   60275 => x"ffffff",
   60276 => x"ffffff",
   60277 => x"ffffff",
   60278 => x"ffffff",
   60279 => x"ffffff",
   60280 => x"ffffff",
   60281 => x"ffffff",
   60282 => x"ffffff",
   60283 => x"ffffff",
   60284 => x"ffffff",
   60285 => x"ffffff",
   60286 => x"ffffff",
   60287 => x"ffffff",
   60288 => x"ffffff",
   60289 => x"ffffff",
   60290 => x"ffffff",
   60291 => x"ffffff",
   60292 => x"ffffff",
   60293 => x"ffffff",
   60294 => x"ffffff",
   60295 => x"ffffff",
   60296 => x"ffffff",
   60297 => x"ffffff",
   60298 => x"ffffff",
   60299 => x"ffffff",
   60300 => x"ffffff",
   60301 => x"ffffff",
   60302 => x"ffffff",
   60303 => x"ffffff",
   60304 => x"ffffff",
   60305 => x"ffffff",
   60306 => x"ffffff",
   60307 => x"ffffff",
   60308 => x"ffffff",
   60309 => x"ffffff",
   60310 => x"ffffff",
   60311 => x"ffffff",
   60312 => x"ffffff",
   60313 => x"ffffff",
   60314 => x"ffffff",
   60315 => x"ffffff",
   60316 => x"ffffff",
   60317 => x"ffffff",
   60318 => x"ffffff",
   60319 => x"ffffff",
   60320 => x"ffffff",
   60321 => x"ffffff",
   60322 => x"ffffff",
   60323 => x"ffffff",
   60324 => x"ffffff",
   60325 => x"ffffff",
   60326 => x"ffffff",
   60327 => x"ffffff",
   60328 => x"ffffff",
   60329 => x"ffffff",
   60330 => x"ffffff",
   60331 => x"ffffff",
   60332 => x"ffffff",
   60333 => x"ffffff",
   60334 => x"ffffff",
   60335 => x"ffffff",
   60336 => x"ffffff",
   60337 => x"ffffff",
   60338 => x"ffffff",
   60339 => x"ffffff",
   60340 => x"ffffff",
   60341 => x"ffffff",
   60342 => x"ffffff",
   60343 => x"ffffff",
   60344 => x"ffffff",
   60345 => x"ffffff",
   60346 => x"ffffff",
   60347 => x"ffffff",
   60348 => x"ffffff",
   60349 => x"ffffff",
   60350 => x"ffffff",
   60351 => x"ffffff",
   60352 => x"ffffff",
   60353 => x"ffffff",
   60354 => x"ffffff",
   60355 => x"ffffff",
   60356 => x"ffffff",
   60357 => x"ffffff",
   60358 => x"ffffff",
   60359 => x"ffffff",
   60360 => x"ffffff",
   60361 => x"ffffff",
   60362 => x"ffffff",
   60363 => x"ffffff",
   60364 => x"ffffff",
   60365 => x"ffffff",
   60366 => x"ffffff",
   60367 => x"ffffff",
   60368 => x"ffffff",
   60369 => x"ffffff",
   60370 => x"ffffff",
   60371 => x"ffffff",
   60372 => x"ffffff",
   60373 => x"ffffff",
   60374 => x"ffffff",
   60375 => x"ffffff",
   60376 => x"ffffff",
   60377 => x"ffffff",
   60378 => x"ffffff",
   60379 => x"ffffff",
   60380 => x"ffffff",
   60381 => x"ffffff",
   60382 => x"ffffff",
   60383 => x"ffffff",
   60384 => x"ffffff",
   60385 => x"ffffff",
   60386 => x"ffffff",
   60387 => x"ffffff",
   60388 => x"ffffff",
   60389 => x"ffffff",
   60390 => x"ffffff",
   60391 => x"ffffff",
   60392 => x"ffffff",
   60393 => x"ffffff",
   60394 => x"ffffff",
   60395 => x"ffffff",
   60396 => x"ffffff",
   60397 => x"ffffff",
   60398 => x"ffffff",
   60399 => x"ffffff",
   60400 => x"ffffff",
   60401 => x"ffffff",
   60402 => x"ffffff",
   60403 => x"ffffff",
   60404 => x"ffffff",
   60405 => x"ffffff",
   60406 => x"ffffff",
   60407 => x"ffffff",
   60408 => x"ffffff",
   60409 => x"ffffff",
   60410 => x"ffffff",
   60411 => x"ffffff",
   60412 => x"ffffff",
   60413 => x"ffffff",
   60414 => x"ffffff",
   60415 => x"ffffff",
   60416 => x"ffffff",
   60417 => x"ffffff",
   60418 => x"ffffff",
   60419 => x"ffffff",
   60420 => x"ffffff",
   60421 => x"ffffff",
   60422 => x"ffffff",
   60423 => x"ffffff",
   60424 => x"ffffff",
   60425 => x"ffffff",
   60426 => x"ffffff",
   60427 => x"ffffff",
   60428 => x"ffffff",
   60429 => x"ffffff",
   60430 => x"ffffff",
   60431 => x"ffffff",
   60432 => x"ffffff",
   60433 => x"ffffff",
   60434 => x"ffffff",
   60435 => x"ffffff",
   60436 => x"ffffff",
   60437 => x"ffffff",
   60438 => x"ffffff",
   60439 => x"ffffff",
   60440 => x"ffffff",
   60441 => x"ffffff",
   60442 => x"ffffff",
   60443 => x"ffffff",
   60444 => x"ffffff",
   60445 => x"ffffff",
   60446 => x"ffffff",
   60447 => x"ffffff",
   60448 => x"ffffff",
   60449 => x"ffffff",
   60450 => x"ffffff",
   60451 => x"ffffff",
   60452 => x"ffffff",
   60453 => x"ffffff",
   60454 => x"ffffff",
   60455 => x"ffffff",
   60456 => x"ffffff",
   60457 => x"ffffff",
   60458 => x"ffffff",
   60459 => x"ffffff",
   60460 => x"ffffff",
   60461 => x"ffffff",
   60462 => x"ffffff",
   60463 => x"ffffff",
   60464 => x"ffffff",
   60465 => x"ffffff",
   60466 => x"ffffff",
   60467 => x"ffffff",
   60468 => x"ffffff",
   60469 => x"ffffff",
   60470 => x"ffffff",
   60471 => x"ffffff",
   60472 => x"ffffff",
   60473 => x"ffffff",
   60474 => x"ffffff",
   60475 => x"ffffff",
   60476 => x"ffffff",
   60477 => x"ffffff",
   60478 => x"ffffff",
   60479 => x"ffffff",
   60480 => x"ffffff",
   60481 => x"ffffff",
   60482 => x"ffffff",
   60483 => x"ffffff",
   60484 => x"ffffff",
   60485 => x"ffffff",
   60486 => x"ffffff",
   60487 => x"ffffff",
   60488 => x"ffffff",
   60489 => x"ffffff",
   60490 => x"ffffff",
   60491 => x"ffffff",
   60492 => x"ffffff",
   60493 => x"ffffff",
   60494 => x"ffffff",
   60495 => x"ffffff",
   60496 => x"ffffff",
   60497 => x"ffffff",
   60498 => x"ffffff",
   60499 => x"ffffff",
   60500 => x"ffffff",
   60501 => x"ffffff",
   60502 => x"ffffff",
   60503 => x"ffffff",
   60504 => x"ffffff",
   60505 => x"ffffff",
   60506 => x"ffffff",
   60507 => x"ffffff",
   60508 => x"ffffff",
   60509 => x"ffffff",
   60510 => x"ffffff",
   60511 => x"ffffff",
   60512 => x"ffffff",
   60513 => x"ffffff",
   60514 => x"ffffff",
   60515 => x"ffffff",
   60516 => x"ffffff",
   60517 => x"ffffff",
   60518 => x"ffffff",
   60519 => x"ffffff",
   60520 => x"ffffff",
   60521 => x"ffffff",
   60522 => x"ffffff",
   60523 => x"ffffff",
   60524 => x"ffffff",
   60525 => x"ffffff",
   60526 => x"ffffff",
   60527 => x"ffffff",
   60528 => x"ffffff",
   60529 => x"ffffff",
   60530 => x"ffffff",
   60531 => x"ffffff",
   60532 => x"ffffff",
   60533 => x"ffffff",
   60534 => x"ffffff",
   60535 => x"ffffff",
   60536 => x"ffffff",
   60537 => x"ffffff",
   60538 => x"ffffff",
   60539 => x"ffffff",
   60540 => x"ffffff",
   60541 => x"ffffff",
   60542 => x"ffffff",
   60543 => x"ffffff",
   60544 => x"ffffff",
   60545 => x"ffffff",
   60546 => x"ffffff",
   60547 => x"ffffff",
   60548 => x"ffffff",
   60549 => x"ffffff",
   60550 => x"ffffff",
   60551 => x"ffffff",
   60552 => x"ffffff",
   60553 => x"ffffff",
   60554 => x"ffffff",
   60555 => x"ffffff",
   60556 => x"ffffff",
   60557 => x"ffffff",
   60558 => x"ffffff",
   60559 => x"ffffff",
   60560 => x"ffffff",
   60561 => x"ffffff",
   60562 => x"ffffff",
   60563 => x"ffffff",
   60564 => x"ffffff",
   60565 => x"ffffff",
   60566 => x"ffffff",
   60567 => x"ffffff",
   60568 => x"ffffff",
   60569 => x"ffffff",
   60570 => x"ffffff",
   60571 => x"ffffff",
   60572 => x"ffffff",
   60573 => x"ffffff",
   60574 => x"ffffff",
   60575 => x"ffffff",
   60576 => x"ffffff",
   60577 => x"ffffff",
   60578 => x"ffffff",
   60579 => x"ffffff",
   60580 => x"ffffff",
   60581 => x"ffffff",
   60582 => x"ffffff",
   60583 => x"ffffff",
   60584 => x"ffffff",
   60585 => x"ffffff",
   60586 => x"ffffff",
   60587 => x"ffffff",
   60588 => x"ffffff",
   60589 => x"ffffff",
   60590 => x"ffffff",
   60591 => x"ffffff",
   60592 => x"ffffff",
   60593 => x"ffffff",
   60594 => x"ffffff",
   60595 => x"ffffff",
   60596 => x"ffffff",
   60597 => x"ffffff",
   60598 => x"ffffff",
   60599 => x"ffffff",
   60600 => x"ffffff",
   60601 => x"ffffff",
   60602 => x"ffffff",
   60603 => x"ffffff",
   60604 => x"ffffff",
   60605 => x"ffffff",
   60606 => x"ffffff",
   60607 => x"ffffff",
   60608 => x"ffffff",
   60609 => x"ffffff",
   60610 => x"ffffff",
   60611 => x"ffffff",
   60612 => x"ffffff",
   60613 => x"ffffff",
   60614 => x"ffffff",
   60615 => x"ffffff",
   60616 => x"ffffff",
   60617 => x"ffffff",
   60618 => x"ffffff",
   60619 => x"ffffff",
   60620 => x"ffffff",
   60621 => x"ffffff",
   60622 => x"ffffff",
   60623 => x"ffffff",
   60624 => x"ffffff",
   60625 => x"ffffff",
   60626 => x"ffffff",
   60627 => x"ffffff",
   60628 => x"ffffff",
   60629 => x"ffffff",
   60630 => x"ffffff",
   60631 => x"ffffff",
   60632 => x"ffffff",
   60633 => x"ffffff",
   60634 => x"ffffff",
   60635 => x"ffffff",
   60636 => x"ffffff",
   60637 => x"ffffff",
   60638 => x"ffffff",
   60639 => x"ffffff",
   60640 => x"ffffff",
   60641 => x"ffffff",
   60642 => x"ffffff",
   60643 => x"ffffff",
   60644 => x"ffffff",
   60645 => x"ffffff",
   60646 => x"ffffff",
   60647 => x"ffffff",
   60648 => x"ffffff",
   60649 => x"ffffff",
   60650 => x"ffffff",
   60651 => x"ffffff",
   60652 => x"ffffff",
   60653 => x"ffffff",
   60654 => x"ffffff",
   60655 => x"ffffff",
   60656 => x"ffffff",
   60657 => x"ffffff",
   60658 => x"ffffff",
   60659 => x"ffffff",
   60660 => x"ffffff",
   60661 => x"ffffff",
   60662 => x"ffffff",
   60663 => x"ffffff",
   60664 => x"ffffff",
   60665 => x"ffffff",
   60666 => x"ffffff",
   60667 => x"ffffff",
   60668 => x"ffffff",
   60669 => x"ffffff",
   60670 => x"ffffff",
   60671 => x"ffffff",
   60672 => x"ffffff",
   60673 => x"ffffff",
   60674 => x"ffffff",
   60675 => x"ffffff",
   60676 => x"ffffff",
   60677 => x"ffffff",
   60678 => x"ffffff",
   60679 => x"ffffff",
   60680 => x"ffffff",
   60681 => x"ffffff",
   60682 => x"ffffff",
   60683 => x"ffffff",
   60684 => x"ffffff",
   60685 => x"ffffff",
   60686 => x"ffffff",
   60687 => x"ffffff",
   60688 => x"ffffff",
   60689 => x"ffffff",
   60690 => x"ffffff",
   60691 => x"ffffff",
   60692 => x"ffffff",
   60693 => x"ffffff",
   60694 => x"ffffff",
   60695 => x"ffffff",
   60696 => x"ffffff",
   60697 => x"ffffff",
   60698 => x"ffffff",
   60699 => x"ffffff",
   60700 => x"ffffff",
   60701 => x"ffffff",
   60702 => x"ffffff",
   60703 => x"ffffff",
   60704 => x"ffffff",
   60705 => x"ffffff",
   60706 => x"ffffff",
   60707 => x"ffffff",
   60708 => x"ffffff",
   60709 => x"ffffff",
   60710 => x"ffffff",
   60711 => x"ffffff",
   60712 => x"ffffff",
   60713 => x"ffffff",
   60714 => x"ffffff",
   60715 => x"ffffff",
   60716 => x"ffffff",
   60717 => x"ffffff",
   60718 => x"ffffff",
   60719 => x"ffffff",
   60720 => x"ffffff",
   60721 => x"ffffff",
   60722 => x"ffffff",
   60723 => x"ffffff",
   60724 => x"ffffff",
   60725 => x"ffffff",
   60726 => x"ffffff",
   60727 => x"ffffff",
   60728 => x"ffffff",
   60729 => x"ffffff",
   60730 => x"ffffff",
   60731 => x"ffffff",
   60732 => x"ffffff",
   60733 => x"ffffff",
   60734 => x"ffffff",
   60735 => x"ffffff",
   60736 => x"ffffff",
   60737 => x"ffffff",
   60738 => x"ffffff",
   60739 => x"ffffff",
   60740 => x"ffffff",
   60741 => x"ffffff",
   60742 => x"ffffff",
   60743 => x"ffffff",
   60744 => x"ffffff",
   60745 => x"ffffff",
   60746 => x"ffffff",
   60747 => x"ffffff",
   60748 => x"ffffff",
   60749 => x"ffffff",
   60750 => x"ffffff",
   60751 => x"ffffff",
   60752 => x"ffffff",
   60753 => x"ffffff",
   60754 => x"ffffff",
   60755 => x"ffffff",
   60756 => x"ffffff",
   60757 => x"ffffff",
   60758 => x"ffffff",
   60759 => x"ffffff",
   60760 => x"ffffff",
   60761 => x"ffffff",
   60762 => x"ffffff",
   60763 => x"ffffff",
   60764 => x"ffffff",
   60765 => x"ffffff",
   60766 => x"ffffff",
   60767 => x"ffffff",
   60768 => x"ffffff",
   60769 => x"ffffff",
   60770 => x"ffffff",
   60771 => x"ffffff",
   60772 => x"ffffff",
   60773 => x"ffffff",
   60774 => x"ffffff",
   60775 => x"ffffff",
   60776 => x"ffffff",
   60777 => x"ffffff",
   60778 => x"ffffff",
   60779 => x"ffffff",
   60780 => x"ffffff",
   60781 => x"ffffff",
   60782 => x"ffffff",
   60783 => x"ffffff",
   60784 => x"ffffff",
   60785 => x"ffffff",
   60786 => x"ffffff",
   60787 => x"ffffff",
   60788 => x"ffffff",
   60789 => x"ffffff",
   60790 => x"ffffff",
   60791 => x"ffffff",
   60792 => x"ffffff",
   60793 => x"ffffff",
   60794 => x"ffffff",
   60795 => x"ffffff",
   60796 => x"ffffff",
   60797 => x"ffffff",
   60798 => x"ffffff",
   60799 => x"ffffff",
   60800 => x"ffffff",
   60801 => x"ffffff",
   60802 => x"ffffff",
   60803 => x"ffffff",
   60804 => x"ffffff",
   60805 => x"ffffff",
   60806 => x"ffffff",
   60807 => x"ffffff",
   60808 => x"ffffff",
   60809 => x"ffffff",
   60810 => x"ffffff",
   60811 => x"ffffff",
   60812 => x"ffffff",
   60813 => x"ffffff",
   60814 => x"ffffff",
   60815 => x"ffffff",
   60816 => x"ffffff",
   60817 => x"ffffff",
   60818 => x"ffffff",
   60819 => x"ffffff",
   60820 => x"ffffff",
   60821 => x"ffffff",
   60822 => x"ffffff",
   60823 => x"ffffff",
   60824 => x"ffffff",
   60825 => x"ffffff",
   60826 => x"ffffff",
   60827 => x"ffffff",
   60828 => x"ffffff",
   60829 => x"ffffff",
   60830 => x"ffffff",
   60831 => x"ffffff",
   60832 => x"ffffff",
   60833 => x"ffffff",
   60834 => x"ffffff",
   60835 => x"ffffff",
   60836 => x"ffffff",
   60837 => x"ffffff",
   60838 => x"ffffff",
   60839 => x"ffffff",
   60840 => x"ffffff",
   60841 => x"ffffff",
   60842 => x"ffffff",
   60843 => x"ffffff",
   60844 => x"ffffff",
   60845 => x"ffffff",
   60846 => x"ffffff",
   60847 => x"ffffff",
   60848 => x"ffffff",
   60849 => x"ffffff",
   60850 => x"ffffff",
   60851 => x"ffffff",
   60852 => x"ffffff",
   60853 => x"ffffff",
   60854 => x"ffffff",
   60855 => x"ffffff",
   60856 => x"ffffff",
   60857 => x"ffffff",
   60858 => x"ffffff",
   60859 => x"ffffff",
   60860 => x"ffffff",
   60861 => x"ffffff",
   60862 => x"ffffff",
   60863 => x"ffffff",
   60864 => x"ffffff",
   60865 => x"ffffff",
   60866 => x"ffffff",
   60867 => x"ffffff",
   60868 => x"ffffff",
   60869 => x"ffffff",
   60870 => x"ffffff",
   60871 => x"ffffff",
   60872 => x"ffffff",
   60873 => x"ffffff",
   60874 => x"ffffff",
   60875 => x"ffffff",
   60876 => x"ffffff",
   60877 => x"ffffff",
   60878 => x"ffffff",
   60879 => x"ffffff",
   60880 => x"ffffff",
   60881 => x"ffffff",
   60882 => x"ffffff",
   60883 => x"ffffff",
   60884 => x"ffffff",
   60885 => x"ffffff",
   60886 => x"ffffff",
   60887 => x"ffffff",
   60888 => x"ffffff",
   60889 => x"ffffff",
   60890 => x"ffffff",
   60891 => x"ffffff",
   60892 => x"ffffff",
   60893 => x"ffffff",
   60894 => x"ffffff",
   60895 => x"ffffff",
   60896 => x"ffffff",
   60897 => x"ffffff",
   60898 => x"ffffff",
   60899 => x"ffffff",
   60900 => x"ffffff",
   60901 => x"ffffff",
   60902 => x"ffffff",
   60903 => x"ffffff",
   60904 => x"ffffff",
   60905 => x"ffffff",
   60906 => x"ffffff",
   60907 => x"ffffff",
   60908 => x"ffffff",
   60909 => x"ffffff",
   60910 => x"ffffff",
   60911 => x"ffffff",
   60912 => x"ffffff",
   60913 => x"ffffff",
   60914 => x"ffffff",
   60915 => x"ffffff",
   60916 => x"ffffff",
   60917 => x"ffffff",
   60918 => x"ffffff",
   60919 => x"ffffff",
   60920 => x"ffffff",
   60921 => x"ffffff",
   60922 => x"ffffff",
   60923 => x"ffffff",
   60924 => x"ffffff",
   60925 => x"ffffff",
   60926 => x"ffffff",
   60927 => x"ffffff",
   60928 => x"ffffff",
   60929 => x"ffffff",
   60930 => x"ffffff",
   60931 => x"ffffff",
   60932 => x"ffffff",
   60933 => x"ffffff",
   60934 => x"ffffff",
   60935 => x"ffffff",
   60936 => x"ffffff",
   60937 => x"ffffff",
   60938 => x"ffffff",
   60939 => x"ffffff",
   60940 => x"ffffff",
   60941 => x"ffffff",
   60942 => x"ffffff",
   60943 => x"ffffff",
   60944 => x"ffffff",
   60945 => x"ffffff",
   60946 => x"ffffff",
   60947 => x"ffffff",
   60948 => x"ffffff",
   60949 => x"ffffff",
   60950 => x"ffffff",
   60951 => x"ffffff",
   60952 => x"ffffff",
   60953 => x"ffffff",
   60954 => x"ffffff",
   60955 => x"ffffff",
   60956 => x"ffffff",
   60957 => x"ffffff",
   60958 => x"ffffff",
   60959 => x"ffffff",
   60960 => x"ffffff",
   60961 => x"ffffff",
   60962 => x"ffffff",
   60963 => x"ffffff",
   60964 => x"ffffff",
   60965 => x"ffffff",
   60966 => x"ffffff",
   60967 => x"ffffff",
   60968 => x"ffffff",
   60969 => x"ffffff",
   60970 => x"ffffff",
   60971 => x"ffffff",
   60972 => x"ffffff",
   60973 => x"ffffff",
   60974 => x"ffffff",
   60975 => x"ffffff",
   60976 => x"ffffff",
   60977 => x"ffffff",
   60978 => x"ffffff",
   60979 => x"ffffff",
   60980 => x"ffffff",
   60981 => x"ffffff",
   60982 => x"ffffff",
   60983 => x"ffffff",
   60984 => x"ffffff",
   60985 => x"ffffff",
   60986 => x"ffffff",
   60987 => x"ffffff",
   60988 => x"ffffff",
   60989 => x"ffffff",
   60990 => x"ffffff",
   60991 => x"ffffff",
   60992 => x"ffffff",
   60993 => x"ffffff",
   60994 => x"ffffff",
   60995 => x"ffffff",
   60996 => x"ffffff",
   60997 => x"ffffff",
   60998 => x"ffffff",
   60999 => x"ffffff",
   61000 => x"ffffff",
   61001 => x"ffffff",
   61002 => x"ffffff",
   61003 => x"ffffff",
   61004 => x"ffffff",
   61005 => x"ffffff",
   61006 => x"ffffff",
   61007 => x"ffffff",
   61008 => x"ffffff",
   61009 => x"ffffff",
   61010 => x"ffffff",
   61011 => x"ffffff",
   61012 => x"ffffff",
   61013 => x"ffffff",
   61014 => x"ffffff",
   61015 => x"ffffff",
   61016 => x"ffffff",
   61017 => x"ffffff",
   61018 => x"ffffff",
   61019 => x"ffffff",
   61020 => x"ffffff",
   61021 => x"ffffff",
   61022 => x"ffffff",
   61023 => x"ffffff",
   61024 => x"ffffff",
   61025 => x"ffffff",
   61026 => x"ffffff",
   61027 => x"ffffff",
   61028 => x"ffffff",
   61029 => x"ffffff",
   61030 => x"ffffff",
   61031 => x"ffffff",
   61032 => x"ffffff",
   61033 => x"ffffff",
   61034 => x"ffffff",
   61035 => x"ffffff",
   61036 => x"ffffff",
   61037 => x"ffffff",
   61038 => x"ffffff",
   61039 => x"ffffff",
   61040 => x"ffffff",
   61041 => x"ffffff",
   61042 => x"ffffff",
   61043 => x"ffffff",
   61044 => x"ffffff",
   61045 => x"ffffff",
   61046 => x"ffffff",
   61047 => x"ffffff",
   61048 => x"ffffff",
   61049 => x"ffffff",
   61050 => x"ffffff",
   61051 => x"ffffff",
   61052 => x"ffffff",
   61053 => x"ffffff",
   61054 => x"ffffff",
   61055 => x"ffffff",
   61056 => x"ffffff",
   61057 => x"ffffff",
   61058 => x"ffffff",
   61059 => x"ffffff",
   61060 => x"ffffff",
   61061 => x"ffffff",
   61062 => x"ffffff",
   61063 => x"ffffff",
   61064 => x"ffffff",
   61065 => x"ffffff",
   61066 => x"ffffff",
   61067 => x"ffffff",
   61068 => x"ffffff",
   61069 => x"ffffff",
   61070 => x"ffffff",
   61071 => x"ffffff",
   61072 => x"ffffff",
   61073 => x"ffffff",
   61074 => x"ffffff",
   61075 => x"ffffff",
   61076 => x"ffffff",
   61077 => x"ffffff",
   61078 => x"ffffff",
   61079 => x"ffffff",
   61080 => x"ffffff",
   61081 => x"ffffff",
   61082 => x"ffffff",
   61083 => x"ffffff",
   61084 => x"ffffff",
   61085 => x"ffffff",
   61086 => x"ffffff",
   61087 => x"ffffff",
   61088 => x"ffffff",
   61089 => x"ffffff",
   61090 => x"ffffff",
   61091 => x"ffffff",
   61092 => x"ffffff",
   61093 => x"ffffff",
   61094 => x"ffffff",
   61095 => x"ffffff",
   61096 => x"ffffff",
   61097 => x"ffffff",
   61098 => x"ffffff",
   61099 => x"ffffff",
   61100 => x"ffffff",
   61101 => x"ffffff",
   61102 => x"ffffff",
   61103 => x"ffffff",
   61104 => x"ffffff",
   61105 => x"ffffff",
   61106 => x"ffffff",
   61107 => x"ffffff",
   61108 => x"ffffff",
   61109 => x"ffffff",
   61110 => x"ffffff",
   61111 => x"ffffff",
   61112 => x"ffffff",
   61113 => x"ffffff",
   61114 => x"ffffff",
   61115 => x"ffffff",
   61116 => x"ffffff",
   61117 => x"ffffff",
   61118 => x"ffffff",
   61119 => x"ffffff",
   61120 => x"ffffff",
   61121 => x"ffffff",
   61122 => x"ffffff",
   61123 => x"ffffff",
   61124 => x"ffffff",
   61125 => x"ffffff",
   61126 => x"ffffff",
   61127 => x"ffffff",
   61128 => x"ffffff",
   61129 => x"ffffff",
   61130 => x"ffffff",
   61131 => x"ffffff",
   61132 => x"ffffff",
   61133 => x"ffffff",
   61134 => x"ffffff",
   61135 => x"ffffff",
   61136 => x"ffffff",
   61137 => x"ffffff",
   61138 => x"ffffff",
   61139 => x"ffffff",
   61140 => x"ffffff",
   61141 => x"ffffff",
   61142 => x"ffffff",
   61143 => x"ffffff",
   61144 => x"ffffff",
   61145 => x"ffffff",
   61146 => x"ffffff",
   61147 => x"ffffff",
   61148 => x"ffffff",
   61149 => x"ffffff",
   61150 => x"ffffff",
   61151 => x"ffffff",
   61152 => x"ffffff",
   61153 => x"ffffff",
   61154 => x"ffffff",
   61155 => x"ffffff",
   61156 => x"ffffff",
   61157 => x"ffffff",
   61158 => x"ffffff",
   61159 => x"ffffff",
   61160 => x"ffffff",
   61161 => x"ffffff",
   61162 => x"ffffff",
   61163 => x"ffffff",
   61164 => x"ffffff",
   61165 => x"ffffff",
   61166 => x"ffffff",
   61167 => x"ffffff",
   61168 => x"ffffff",
   61169 => x"ffffff",
   61170 => x"ffffff",
   61171 => x"ffffff",
   61172 => x"ffffff",
   61173 => x"ffffff",
   61174 => x"ffffff",
   61175 => x"ffffff",
   61176 => x"ffffff",
   61177 => x"ffffff",
   61178 => x"ffffff",
   61179 => x"ffffff",
   61180 => x"ffffff",
   61181 => x"ffffff",
   61182 => x"ffffff",
   61183 => x"ffffff",
   61184 => x"ffffff",
   61185 => x"ffffff",
   61186 => x"ffffff",
   61187 => x"ffffff",
   61188 => x"ffffff",
   61189 => x"ffffff",
   61190 => x"ffffff",
   61191 => x"ffffff",
   61192 => x"ffffff",
   61193 => x"ffffff",
   61194 => x"ffffff",
   61195 => x"ffffff",
   61196 => x"ffffff",
   61197 => x"ffffff",
   61198 => x"ffffff",
   61199 => x"ffffff",
   61200 => x"ffffff",
   61201 => x"ffffff",
   61202 => x"ffffff",
   61203 => x"ffffff",
   61204 => x"ffffff",
   61205 => x"ffffff",
   61206 => x"ffffff",
   61207 => x"ffffff",
   61208 => x"ffffff",
   61209 => x"ffffff",
   61210 => x"ffffff",
   61211 => x"ffffff",
   61212 => x"ffffff",
   61213 => x"ffffff",
   61214 => x"ffffff",
   61215 => x"ffffff",
   61216 => x"ffffff",
   61217 => x"ffffff",
   61218 => x"ffffff",
   61219 => x"ffffff",
   61220 => x"ffffff",
   61221 => x"ffffff",
   61222 => x"ffffff",
   61223 => x"ffffff",
   61224 => x"ffffff",
   61225 => x"ffffff",
   61226 => x"ffffff",
   61227 => x"ffffff",
   61228 => x"ffffff",
   61229 => x"ffffff",
   61230 => x"ffffff",
   61231 => x"ffffff",
   61232 => x"ffffff",
   61233 => x"ffffff",
   61234 => x"ffffff",
   61235 => x"ffffff",
   61236 => x"ffffff",
   61237 => x"ffffff",
   61238 => x"ffffff",
   61239 => x"ffffff",
   61240 => x"ffffff",
   61241 => x"ffffff",
   61242 => x"ffffff",
   61243 => x"ffffff",
   61244 => x"ffffff",
   61245 => x"ffffff",
   61246 => x"ffffff",
   61247 => x"ffffff",
   61248 => x"ffffff",
   61249 => x"ffffff",
   61250 => x"ffffff",
   61251 => x"ffffff",
   61252 => x"ffffff",
   61253 => x"ffffff",
   61254 => x"ffffff",
   61255 => x"ffffff",
   61256 => x"ffffff",
   61257 => x"ffffff",
   61258 => x"ffffff",
   61259 => x"ffffff",
   61260 => x"ffffff",
   61261 => x"ffffff",
   61262 => x"ffffff",
   61263 => x"ffffff",
   61264 => x"ffffff",
   61265 => x"ffffff",
   61266 => x"ffffff",
   61267 => x"ffffff",
   61268 => x"ffffff",
   61269 => x"ffffff",
   61270 => x"ffffff",
   61271 => x"ffffff",
   61272 => x"ffffff",
   61273 => x"ffffff",
   61274 => x"ffffff",
   61275 => x"ffffff",
   61276 => x"ffffff",
   61277 => x"ffffff",
   61278 => x"ffffff",
   61279 => x"ffffff",
   61280 => x"ffffff",
   61281 => x"ffffff",
   61282 => x"ffffff",
   61283 => x"ffffff",
   61284 => x"ffffff",
   61285 => x"ffffff",
   61286 => x"ffffff",
   61287 => x"ffffff",
   61288 => x"ffffff",
   61289 => x"ffffff",
   61290 => x"ffffff",
   61291 => x"ffffff",
   61292 => x"ffffff",
   61293 => x"ffffff",
   61294 => x"ffffff",
   61295 => x"ffffff",
   61296 => x"ffffff",
   61297 => x"ffffff",
   61298 => x"ffffff",
   61299 => x"ffffff",
   61300 => x"ffffff",
   61301 => x"ffffff",
   61302 => x"ffffff",
   61303 => x"ffffff",
   61304 => x"ffffff",
   61305 => x"ffffff",
   61306 => x"ffffff",
   61307 => x"ffffff",
   61308 => x"ffffff",
   61309 => x"ffffff",
   61310 => x"ffffff",
   61311 => x"ffffff",
   61312 => x"ffffff",
   61313 => x"ffffff",
   61314 => x"ffffff",
   61315 => x"ffffff",
   61316 => x"ffffff",
   61317 => x"ffffff",
   61318 => x"ffffff",
   61319 => x"ffffff",
   61320 => x"ffffff",
   61321 => x"ffffff",
   61322 => x"ffffff",
   61323 => x"ffffff",
   61324 => x"ffffff",
   61325 => x"ffffff",
   61326 => x"ffffff",
   61327 => x"ffffff",
   61328 => x"ffffff",
   61329 => x"ffffff",
   61330 => x"ffffff",
   61331 => x"ffffff",
   61332 => x"ffffff",
   61333 => x"ffffff",
   61334 => x"ffffff",
   61335 => x"ffffff",
   61336 => x"ffffff",
   61337 => x"ffffff",
   61338 => x"ffffff",
   61339 => x"ffffff",
   61340 => x"ffffff",
   61341 => x"ffffff",
   61342 => x"ffffff",
   61343 => x"ffffff",
   61344 => x"ffffff",
   61345 => x"ffffff",
   61346 => x"ffffff",
   61347 => x"ffffff",
   61348 => x"ffffff",
   61349 => x"ffffff",
   61350 => x"ffffff",
   61351 => x"ffffff",
   61352 => x"ffffff",
   61353 => x"ffffff",
   61354 => x"ffffff",
   61355 => x"ffffff",
   61356 => x"ffffff",
   61357 => x"ffffff",
   61358 => x"ffffff",
   61359 => x"ffffff",
   61360 => x"ffffff",
   61361 => x"ffffff",
   61362 => x"ffffff",
   61363 => x"ffffff",
   61364 => x"ffffff",
   61365 => x"ffffff",
   61366 => x"ffffff",
   61367 => x"ffffff",
   61368 => x"ffffff",
   61369 => x"ffffff",
   61370 => x"ffffff",
   61371 => x"ffffff",
   61372 => x"ffffff",
   61373 => x"ffffff",
   61374 => x"ffffff",
   61375 => x"ffffff",
   61376 => x"ffffff",
   61377 => x"ffffff",
   61378 => x"ffffff",
   61379 => x"ffffff",
   61380 => x"ffffff",
   61381 => x"ffffff",
   61382 => x"ffffff",
   61383 => x"ffffff",
   61384 => x"ffffff",
   61385 => x"ffffff",
   61386 => x"ffffff",
   61387 => x"ffffff",
   61388 => x"ffffff",
   61389 => x"ffffff",
   61390 => x"ffffff",
   61391 => x"ffffff",
   61392 => x"ffffff",
   61393 => x"ffffff",
   61394 => x"ffffff",
   61395 => x"ffffff",
   61396 => x"ffffff",
   61397 => x"ffffff",
   61398 => x"ffffff",
   61399 => x"ffffff",
   61400 => x"ffffff",
   61401 => x"ffffff",
   61402 => x"ffffff",
   61403 => x"ffffff",
   61404 => x"ffffff",
   61405 => x"ffffff",
   61406 => x"ffffff",
   61407 => x"ffffff",
   61408 => x"ffffff",
   61409 => x"ffffff",
   61410 => x"ffffff",
   61411 => x"ffffff",
   61412 => x"ffffff",
   61413 => x"ffffff",
   61414 => x"ffffff",
   61415 => x"ffffff",
   61416 => x"ffffff",
   61417 => x"ffffff",
   61418 => x"ffffff",
   61419 => x"ffffff",
   61420 => x"ffffff",
   61421 => x"ffffff",
   61422 => x"ffffff",
   61423 => x"ffffff",
   61424 => x"ffffff",
   61425 => x"ffffff",
   61426 => x"ffffff",
   61427 => x"ffffff",
   61428 => x"ffffff",
   61429 => x"ffffff",
   61430 => x"ffffff",
   61431 => x"ffffff",
   61432 => x"ffffff",
   61433 => x"ffffff",
   61434 => x"ffffff",
   61435 => x"ffffff",
   61436 => x"ffffff",
   61437 => x"ffffff",
   61438 => x"ffffff",
   61439 => x"ffffff",
   61440 => x"ffffff",
   61441 => x"ffffff",
   61442 => x"ffffff",
   61443 => x"ffffff",
   61444 => x"ffffff",
   61445 => x"ffffff",
   61446 => x"ffffff",
   61447 => x"ffffff",
   61448 => x"ffffff",
   61449 => x"ffffff",
   61450 => x"ffffff",
   61451 => x"ffffff",
   61452 => x"ffffff",
   61453 => x"ffffff",
   61454 => x"ffffff",
   61455 => x"ffffff",
   61456 => x"ffffff",
   61457 => x"ffffff",
   61458 => x"ffffff",
   61459 => x"ffffff",
   61460 => x"ffffff",
   61461 => x"ffffff",
   61462 => x"ffffff",
   61463 => x"ffffff",
   61464 => x"ffffff",
   61465 => x"ffffff",
   61466 => x"ffffff",
   61467 => x"ffffff",
   61468 => x"ffffff",
   61469 => x"ffffff",
   61470 => x"ffffff",
   61471 => x"ffffff",
   61472 => x"ffffff",
   61473 => x"ffffff",
   61474 => x"ffffff",
   61475 => x"ffffff",
   61476 => x"ffffff",
   61477 => x"ffffff",
   61478 => x"ffffff",
   61479 => x"ffffff",
   61480 => x"ffffff",
   61481 => x"ffffff",
   61482 => x"ffffff",
   61483 => x"ffffff",
   61484 => x"ffffff",
   61485 => x"ffffff",
   61486 => x"ffffff",
   61487 => x"ffffff",
   61488 => x"ffffff",
   61489 => x"ffffff",
   61490 => x"ffffff",
   61491 => x"ffffff",
   61492 => x"ffffff",
   61493 => x"ffffff",
   61494 => x"ffffff",
   61495 => x"ffffff",
   61496 => x"ffffff",
   61497 => x"ffffff",
   61498 => x"ffffff",
   61499 => x"ffffff",
   61500 => x"ffffff",
   61501 => x"ffffff",
   61502 => x"ffffff",
   61503 => x"ffffff",
   61504 => x"ffffff",
   61505 => x"ffffff",
   61506 => x"ffffff",
   61507 => x"ffffff",
   61508 => x"ffffff",
   61509 => x"ffffff",
   61510 => x"ffffff",
   61511 => x"ffffff",
   61512 => x"ffffff",
   61513 => x"ffffff",
   61514 => x"ffffff",
   61515 => x"ffffff",
   61516 => x"ffffff",
   61517 => x"ffffff",
   61518 => x"ffffff",
   61519 => x"ffffff",
   61520 => x"ffffff",
   61521 => x"ffffff",
   61522 => x"ffffff",
   61523 => x"ffffff",
   61524 => x"ffffff",
   61525 => x"ffffff",
   61526 => x"ffffff",
   61527 => x"ffffff",
   61528 => x"ffffff",
   61529 => x"ffffff",
   61530 => x"ffffff",
   61531 => x"ffffff",
   61532 => x"ffffff",
   61533 => x"ffffff",
   61534 => x"ffffff",
   61535 => x"ffffff",
   61536 => x"ffffff",
   61537 => x"ffffff",
   61538 => x"ffffff",
   61539 => x"ffffff",
   61540 => x"ffffff",
   61541 => x"ffffff",
   61542 => x"ffffff",
   61543 => x"ffffff",
   61544 => x"ffffff",
   61545 => x"ffffff",
   61546 => x"ffffff",
   61547 => x"ffffff",
   61548 => x"ffffff",
   61549 => x"ffffff",
   61550 => x"ffffff",
   61551 => x"ffffff",
   61552 => x"ffffff",
   61553 => x"ffffff",
   61554 => x"ffffff",
   61555 => x"ffffff",
   61556 => x"ffffff",
   61557 => x"ffffff",
   61558 => x"ffffff",
   61559 => x"ffffff",
   61560 => x"ffffff",
   61561 => x"ffffff",
   61562 => x"ffffff",
   61563 => x"ffffff",
   61564 => x"ffffff",
   61565 => x"ffffff",
   61566 => x"ffffff",
   61567 => x"ffffff",
   61568 => x"ffffff",
   61569 => x"ffffff",
   61570 => x"ffffff",
   61571 => x"ffffff",
   61572 => x"ffffff",
   61573 => x"ffffff",
   61574 => x"ffffff",
   61575 => x"ffffff",
   61576 => x"ffffff",
   61577 => x"ffffff",
   61578 => x"ffffff",
   61579 => x"ffffff",
   61580 => x"ffffff",
   61581 => x"ffffff",
   61582 => x"ffffff",
   61583 => x"ffffff",
   61584 => x"ffffff",
   61585 => x"ffffff",
   61586 => x"ffffff",
   61587 => x"ffffff",
   61588 => x"ffffff",
   61589 => x"ffffff",
   61590 => x"ffffff",
   61591 => x"ffffff",
   61592 => x"ffffff",
   61593 => x"ffffff",
   61594 => x"ffffff",
   61595 => x"ffffff",
   61596 => x"ffffff",
   61597 => x"ffffff",
   61598 => x"ffffff",
   61599 => x"ffffff",
   61600 => x"ffffff",
   61601 => x"ffffff",
   61602 => x"ffffff",
   61603 => x"ffffff",
   61604 => x"ffffff",
   61605 => x"ffffff",
   61606 => x"ffffff",
   61607 => x"ffffff",
   61608 => x"ffffff",
   61609 => x"ffffff",
   61610 => x"ffffff",
   61611 => x"ffffff",
   61612 => x"ffffff",
   61613 => x"ffffff",
   61614 => x"ffffff",
   61615 => x"ffffff",
   61616 => x"ffffff",
   61617 => x"ffffff",
   61618 => x"ffffff",
   61619 => x"ffffff",
   61620 => x"ffffff",
   61621 => x"ffffff",
   61622 => x"ffffff",
   61623 => x"ffffff",
   61624 => x"ffffff",
   61625 => x"ffffff",
   61626 => x"ffffff",
   61627 => x"ffffff",
   61628 => x"ffffff",
   61629 => x"ffffff",
   61630 => x"ffffff",
   61631 => x"ffffff",
   61632 => x"ffffff",
   61633 => x"ffffff",
   61634 => x"ffffff",
   61635 => x"ffffff",
   61636 => x"ffffff",
   61637 => x"ffffff",
   61638 => x"ffffff",
   61639 => x"ffffff",
   61640 => x"ffffff",
   61641 => x"ffffff",
   61642 => x"ffffff",
   61643 => x"ffffff",
   61644 => x"ffffff",
   61645 => x"ffffff",
   61646 => x"ffffff",
   61647 => x"ffffff",
   61648 => x"ffffff",
   61649 => x"ffffff",
   61650 => x"ffffff",
   61651 => x"ffffff",
   61652 => x"ffffff",
   61653 => x"ffffff",
   61654 => x"ffffff",
   61655 => x"ffffff",
   61656 => x"ffffff",
   61657 => x"ffffff",
   61658 => x"ffffff",
   61659 => x"ffffff",
   61660 => x"ffffff",
   61661 => x"ffffff",
   61662 => x"ffffff",
   61663 => x"ffffff",
   61664 => x"ffffff",
   61665 => x"ffffff",
   61666 => x"ffffff",
   61667 => x"ffffff",
   61668 => x"ffffff",
   61669 => x"ffffff",
   61670 => x"ffffff",
   61671 => x"ffffff",
   61672 => x"ffffff",
   61673 => x"ffffff",
   61674 => x"ffffff",
   61675 => x"ffffff",
   61676 => x"ffffff",
   61677 => x"ffffff",
   61678 => x"ffffff",
   61679 => x"ffffff",
   61680 => x"ffffff",
   61681 => x"ffffff",
   61682 => x"ffffff",
   61683 => x"ffffff",
   61684 => x"ffffff",
   61685 => x"ffffff",
   61686 => x"ffffff",
   61687 => x"ffffff",
   61688 => x"ffffff",
   61689 => x"ffffff",
   61690 => x"ffffff",
   61691 => x"ffffff",
   61692 => x"ffffff",
   61693 => x"ffffff",
   61694 => x"ffffff",
   61695 => x"ffffff",
   61696 => x"ffffff",
   61697 => x"ffffff",
   61698 => x"ffffff",
   61699 => x"ffffff",
   61700 => x"ffffff",
   61701 => x"ffffff",
   61702 => x"ffffff",
   61703 => x"ffffff",
   61704 => x"ffffff",
   61705 => x"ffffff",
   61706 => x"ffffff",
   61707 => x"ffffff",
   61708 => x"ffffff",
   61709 => x"ffffff",
   61710 => x"ffffff",
   61711 => x"ffffff",
   61712 => x"ffffff",
   61713 => x"ffffff",
   61714 => x"ffffff",
   61715 => x"ffffff",
   61716 => x"ffffff",
   61717 => x"ffffff",
   61718 => x"ffffff",
   61719 => x"ffffff",
   61720 => x"ffffff",
   61721 => x"ffffff",
   61722 => x"ffffff",
   61723 => x"ffffff",
   61724 => x"ffffff",
   61725 => x"ffffff",
   61726 => x"ffffff",
   61727 => x"ffffff",
   61728 => x"ffffff",
   61729 => x"ffffff",
   61730 => x"ffffff",
   61731 => x"ffffff",
   61732 => x"ffffff",
   61733 => x"ffffff",
   61734 => x"ffffff",
   61735 => x"ffffff",
   61736 => x"ffffff",
   61737 => x"ffffff",
   61738 => x"ffffff",
   61739 => x"ffffff",
   61740 => x"ffffff",
   61741 => x"ffffff",
   61742 => x"ffffff",
   61743 => x"ffffff",
   61744 => x"ffffff",
   61745 => x"ffffff",
   61746 => x"ffffff",
   61747 => x"ffffff",
   61748 => x"ffffff",
   61749 => x"ffffff",
   61750 => x"ffffff",
   61751 => x"ffffff",
   61752 => x"ffffff",
   61753 => x"ffffff",
   61754 => x"ffffff",
   61755 => x"ffffff",
   61756 => x"ffffff",
   61757 => x"ffffff",
   61758 => x"ffffff",
   61759 => x"ffffff",
   61760 => x"ffffff",
   61761 => x"ffffff",
   61762 => x"ffffff",
   61763 => x"ffffff",
   61764 => x"ffffff",
   61765 => x"ffffff",
   61766 => x"ffffff",
   61767 => x"ffffff",
   61768 => x"ffffff",
   61769 => x"ffffff",
   61770 => x"ffffff",
   61771 => x"ffffff",
   61772 => x"ffffff",
   61773 => x"ffffff",
   61774 => x"ffffff",
   61775 => x"ffffff",
   61776 => x"ffffff",
   61777 => x"ffffff",
   61778 => x"ffffff",
   61779 => x"ffffff",
   61780 => x"ffffff",
   61781 => x"ffffff",
   61782 => x"ffffff",
   61783 => x"ffffff",
   61784 => x"ffffff",
   61785 => x"ffffff",
   61786 => x"ffffff",
   61787 => x"ffffff",
   61788 => x"ffffff",
   61789 => x"ffffff",
   61790 => x"ffffff",
   61791 => x"ffffff",
   61792 => x"ffffff",
   61793 => x"ffffff",
   61794 => x"ffffff",
   61795 => x"ffffff",
   61796 => x"ffffff",
   61797 => x"ffffff",
   61798 => x"ffffff",
   61799 => x"ffffff",
   61800 => x"ffffff",
   61801 => x"ffffff",
   61802 => x"ffffff",
   61803 => x"ffffff",
   61804 => x"ffffff",
   61805 => x"ffffff",
   61806 => x"ffffff",
   61807 => x"ffffff",
   61808 => x"ffffff",
   61809 => x"ffffff",
   61810 => x"ffffff",
   61811 => x"ffffff",
   61812 => x"ffffff",
   61813 => x"ffffff",
   61814 => x"ffffff",
   61815 => x"ffffff",
   61816 => x"ffffff",
   61817 => x"ffffff",
   61818 => x"ffffff",
   61819 => x"ffffff",
   61820 => x"ffffff",
   61821 => x"ffffff",
   61822 => x"ffffff",
   61823 => x"ffffff",
   61824 => x"ffffff",
   61825 => x"ffffff",
   61826 => x"ffffff",
   61827 => x"ffffff",
   61828 => x"ffffff",
   61829 => x"ffffff",
   61830 => x"ffffff",
   61831 => x"ffffff",
   61832 => x"ffffff",
   61833 => x"ffffff",
   61834 => x"ffffff",
   61835 => x"ffffff",
   61836 => x"ffffff",
   61837 => x"ffffff",
   61838 => x"ffffff",
   61839 => x"ffffff",
   61840 => x"ffffff",
   61841 => x"ffffff",
   61842 => x"ffffff",
   61843 => x"ffffff",
   61844 => x"ffffff",
   61845 => x"ffffff",
   61846 => x"ffffff",
   61847 => x"ffffff",
   61848 => x"ffffff",
   61849 => x"ffffff",
   61850 => x"ffffff",
   61851 => x"ffffff",
   61852 => x"ffffff",
   61853 => x"ffffff",
   61854 => x"ffffff",
   61855 => x"ffffff",
   61856 => x"ffffff",
   61857 => x"ffffff",
   61858 => x"ffffff",
   61859 => x"ffffff",
   61860 => x"ffffff",
   61861 => x"ffffff",
   61862 => x"ffffff",
   61863 => x"ffffff",
   61864 => x"ffffff",
   61865 => x"ffffff",
   61866 => x"ffffff",
   61867 => x"ffffff",
   61868 => x"ffffff",
   61869 => x"ffffff",
   61870 => x"ffffff",
   61871 => x"ffffff",
   61872 => x"ffffff",
   61873 => x"ffffff",
   61874 => x"ffffff",
   61875 => x"ffffff",
   61876 => x"ffffff",
   61877 => x"ffffff",
   61878 => x"ffffff",
   61879 => x"ffffff",
   61880 => x"ffffff",
   61881 => x"ffffff",
   61882 => x"ffffff",
   61883 => x"ffffff",
   61884 => x"ffffff",
   61885 => x"ffffff",
   61886 => x"ffffff",
   61887 => x"ffffff",
   61888 => x"ffffff",
   61889 => x"ffffff",
   61890 => x"ffffff",
   61891 => x"ffffff",
   61892 => x"ffffff",
   61893 => x"ffffff",
   61894 => x"ffffff",
   61895 => x"ffffff",
   61896 => x"ffffff",
   61897 => x"ffffff",
   61898 => x"ffffff",
   61899 => x"ffffff",
   61900 => x"ffffff",
   61901 => x"ffffff",
   61902 => x"ffffff",
   61903 => x"ffffff",
   61904 => x"ffffff",
   61905 => x"ffffff",
   61906 => x"ffffff",
   61907 => x"ffffff",
   61908 => x"ffffff",
   61909 => x"ffffff",
   61910 => x"ffffff",
   61911 => x"ffffff",
   61912 => x"ffffff",
   61913 => x"ffffff",
   61914 => x"ffffff",
   61915 => x"ffffff",
   61916 => x"ffffff",
   61917 => x"ffffff",
   61918 => x"ffffff",
   61919 => x"ffffff",
   61920 => x"ffffff",
   61921 => x"ffffff",
   61922 => x"ffffff",
   61923 => x"ffffff",
   61924 => x"ffffff",
   61925 => x"ffffff",
   61926 => x"ffffff",
   61927 => x"ffffff",
   61928 => x"ffffff",
   61929 => x"ffffff",
   61930 => x"ffffff",
   61931 => x"ffffff",
   61932 => x"ffffff",
   61933 => x"ffffff",
   61934 => x"ffffff",
   61935 => x"ffffff",
   61936 => x"ffffff",
   61937 => x"ffffff",
   61938 => x"ffffff",
   61939 => x"ffffff",
   61940 => x"ffffff",
   61941 => x"ffffff",
   61942 => x"ffffff",
   61943 => x"ffffff",
   61944 => x"ffffff",
   61945 => x"ffffff",
   61946 => x"ffffff",
   61947 => x"ffffff",
   61948 => x"ffffff",
   61949 => x"ffffff",
   61950 => x"ffffff",
   61951 => x"ffffff",
   61952 => x"ffffff",
   61953 => x"ffffff",
   61954 => x"ffffff",
   61955 => x"ffffff",
   61956 => x"ffffff",
   61957 => x"ffffff",
   61958 => x"ffffff",
   61959 => x"ffffff",
   61960 => x"ffffff",
   61961 => x"ffffff",
   61962 => x"ffffff",
   61963 => x"ffffff",
   61964 => x"ffffff",
   61965 => x"ffffff",
   61966 => x"ffffff",
   61967 => x"ffffff",
   61968 => x"ffffff",
   61969 => x"ffffff",
   61970 => x"ffffff",
   61971 => x"ffffff",
   61972 => x"ffffff",
   61973 => x"ffffff",
   61974 => x"ffffff",
   61975 => x"ffffff",
   61976 => x"ffffff",
   61977 => x"ffffff",
   61978 => x"ffffff",
   61979 => x"ffffff",
   61980 => x"ffffff",
   61981 => x"ffffff",
   61982 => x"ffffff",
   61983 => x"ffffff",
   61984 => x"ffffff",
   61985 => x"ffffff",
   61986 => x"ffffff",
   61987 => x"ffffff",
   61988 => x"ffffff",
   61989 => x"ffffff",
   61990 => x"ffffff",
   61991 => x"ffffff",
   61992 => x"ffffff",
   61993 => x"ffffff",
   61994 => x"ffffff",
   61995 => x"ffffff",
   61996 => x"ffffff",
   61997 => x"ffffff",
   61998 => x"ffffff",
   61999 => x"ffffff",
   62000 => x"ffffff",
   62001 => x"ffffff",
   62002 => x"ffffff",
   62003 => x"ffffff",
   62004 => x"ffffff",
   62005 => x"ffffff",
   62006 => x"ffffff",
   62007 => x"ffffff",
   62008 => x"ffffff",
   62009 => x"ffffff",
   62010 => x"ffffff",
   62011 => x"ffffff",
   62012 => x"ffffff",
   62013 => x"ffffff",
   62014 => x"ffffff",
   62015 => x"ffffff",
   62016 => x"ffffff",
   62017 => x"ffffff",
   62018 => x"ffffff",
   62019 => x"ffffff",
   62020 => x"ffffff",
   62021 => x"ffffff",
   62022 => x"ffffff",
   62023 => x"ffffff",
   62024 => x"ffffff",
   62025 => x"ffffff",
   62026 => x"ffffff",
   62027 => x"ffffff",
   62028 => x"ffffff",
   62029 => x"ffffff",
   62030 => x"ffffff",
   62031 => x"ffffff",
   62032 => x"ffffff",
   62033 => x"ffffff",
   62034 => x"ffffff",
   62035 => x"ffffff",
   62036 => x"ffffff",
   62037 => x"ffffff",
   62038 => x"ffffff",
   62039 => x"ffffff",
   62040 => x"ffffff",
   62041 => x"ffffff",
   62042 => x"ffffff",
   62043 => x"ffffff",
   62044 => x"ffffff",
   62045 => x"ffffff",
   62046 => x"ffffff",
   62047 => x"ffffff",
   62048 => x"ffffff",
   62049 => x"ffffff",
   62050 => x"ffffff",
   62051 => x"ffffff",
   62052 => x"ffffff",
   62053 => x"ffffff",
   62054 => x"ffffff",
   62055 => x"ffffff",
   62056 => x"ffffff",
   62057 => x"ffffff",
   62058 => x"ffffff",
   62059 => x"ffffff",
   62060 => x"ffffff",
   62061 => x"ffffff",
   62062 => x"ffffff",
   62063 => x"ffffff",
   62064 => x"ffffff",
   62065 => x"ffffff",
   62066 => x"ffffff",
   62067 => x"ffffff",
   62068 => x"ffffff",
   62069 => x"ffffff",
   62070 => x"ffffff",
   62071 => x"ffffff",
   62072 => x"ffffff",
   62073 => x"ffffff",
   62074 => x"ffffff",
   62075 => x"ffffff",
   62076 => x"ffffff",
   62077 => x"ffffff",
   62078 => x"ffffff",
   62079 => x"ffffff",
   62080 => x"ffffff",
   62081 => x"ffffff",
   62082 => x"ffffff",
   62083 => x"ffffff",
   62084 => x"ffffff",
   62085 => x"ffffff",
   62086 => x"ffffff",
   62087 => x"ffffff",
   62088 => x"ffffff",
   62089 => x"ffffff",
   62090 => x"ffffff",
   62091 => x"ffffff",
   62092 => x"ffffff",
   62093 => x"ffffff",
   62094 => x"ffffff",
   62095 => x"ffffff",
   62096 => x"ffffff",
   62097 => x"ffffff",
   62098 => x"ffffff",
   62099 => x"ffffff",
   62100 => x"ffffff",
   62101 => x"ffffff",
   62102 => x"ffffff",
   62103 => x"ffffff",
   62104 => x"ffffff",
   62105 => x"ffffff",
   62106 => x"ffffff",
   62107 => x"ffffff",
   62108 => x"ffffff",
   62109 => x"ffffff",
   62110 => x"ffffff",
   62111 => x"ffffff",
   62112 => x"ffffff",
   62113 => x"ffffff",
   62114 => x"ffffff",
   62115 => x"ffffff",
   62116 => x"ffffff",
   62117 => x"ffffff",
   62118 => x"ffffff",
   62119 => x"ffffff",
   62120 => x"ffffff",
   62121 => x"ffffff",
   62122 => x"ffffff",
   62123 => x"ffffff",
   62124 => x"ffffff",
   62125 => x"ffffff",
   62126 => x"ffffff",
   62127 => x"ffffff",
   62128 => x"ffffff",
   62129 => x"ffffff",
   62130 => x"ffffff",
   62131 => x"ffffff",
   62132 => x"ffffff",
   62133 => x"ffffff",
   62134 => x"ffffff",
   62135 => x"ffffff",
   62136 => x"ffffff",
   62137 => x"ffffff",
   62138 => x"ffffff",
   62139 => x"ffffff",
   62140 => x"ffffff",
   62141 => x"ffffff",
   62142 => x"ffffff",
   62143 => x"ffffff",
   62144 => x"ffffff",
   62145 => x"ffffff",
   62146 => x"ffffff",
   62147 => x"ffffff",
   62148 => x"ffffff",
   62149 => x"ffffff",
   62150 => x"ffffff",
   62151 => x"ffffff",
   62152 => x"ffffff",
   62153 => x"ffffff",
   62154 => x"ffffff",
   62155 => x"ffffff",
   62156 => x"ffffff",
   62157 => x"ffffff",
   62158 => x"ffffff",
   62159 => x"ffffff",
   62160 => x"ffffff",
   62161 => x"ffffff",
   62162 => x"ffffff",
   62163 => x"ffffff",
   62164 => x"ffffff",
   62165 => x"ffffff",
   62166 => x"ffffff",
   62167 => x"ffffff",
   62168 => x"ffffff",
   62169 => x"ffffff",
   62170 => x"ffffff",
   62171 => x"ffffff",
   62172 => x"ffffff",
   62173 => x"ffffff",
   62174 => x"ffffff",
   62175 => x"ffffff",
   62176 => x"ffffff",
   62177 => x"ffffff",
   62178 => x"ffffff",
   62179 => x"ffffff",
   62180 => x"ffffff",
   62181 => x"ffffff",
   62182 => x"ffffff",
   62183 => x"ffffff",
   62184 => x"ffffff",
   62185 => x"ffffff",
   62186 => x"ffffff",
   62187 => x"ffffff",
   62188 => x"ffffff",
   62189 => x"ffffff",
   62190 => x"ffffff",
   62191 => x"ffffff",
   62192 => x"ffffff",
   62193 => x"ffffff",
   62194 => x"ffffff",
   62195 => x"ffffff",
   62196 => x"ffffff",
   62197 => x"ffffff",
   62198 => x"ffffff",
   62199 => x"ffffff",
   62200 => x"ffffff",
   62201 => x"ffffff",
   62202 => x"ffffff",
   62203 => x"ffffff",
   62204 => x"ffffff",
   62205 => x"ffffff",
   62206 => x"ffffff",
   62207 => x"ffffff",
   62208 => x"ffffff",
   62209 => x"ffffff",
   62210 => x"ffffff",
   62211 => x"ffffff",
   62212 => x"ffffff",
   62213 => x"ffffff",
   62214 => x"ffffff",
   62215 => x"ffffff",
   62216 => x"ffffff",
   62217 => x"ffffff",
   62218 => x"ffffff",
   62219 => x"ffffff",
   62220 => x"ffffff",
   62221 => x"ffffff",
   62222 => x"ffffff",
   62223 => x"ffffff",
   62224 => x"ffffff",
   62225 => x"ffffff",
   62226 => x"ffffff",
   62227 => x"ffffff",
   62228 => x"ffffff",
   62229 => x"ffffff",
   62230 => x"ffffff",
   62231 => x"ffffff",
   62232 => x"ffffff",
   62233 => x"ffffff",
   62234 => x"ffffff",
   62235 => x"ffffff",
   62236 => x"ffffff",
   62237 => x"ffffff",
   62238 => x"ffffff",
   62239 => x"ffffff",
   62240 => x"ffffff",
   62241 => x"ffffff",
   62242 => x"ffffff",
   62243 => x"ffffff",
   62244 => x"ffffff",
   62245 => x"ffffff",
   62246 => x"ffffff",
   62247 => x"ffffff",
   62248 => x"ffffff",
   62249 => x"ffffff",
   62250 => x"ffffff",
   62251 => x"ffffff",
   62252 => x"ffffff",
   62253 => x"ffffff",
   62254 => x"ffffff",
   62255 => x"ffffff",
   62256 => x"ffffff",
   62257 => x"ffffff",
   62258 => x"ffffff",
   62259 => x"ffffff",
   62260 => x"ffffff",
   62261 => x"ffffff",
   62262 => x"ffffff",
   62263 => x"ffffff",
   62264 => x"ffffff",
   62265 => x"ffffff",
   62266 => x"ffffff",
   62267 => x"ffffff",
   62268 => x"ffffff",
   62269 => x"ffffff",
   62270 => x"ffffff",
   62271 => x"ffffff",
   62272 => x"ffffff",
   62273 => x"ffffff",
   62274 => x"ffffff",
   62275 => x"ffffff",
   62276 => x"ffffff",
   62277 => x"ffffff",
   62278 => x"ffffff",
   62279 => x"ffffff",
   62280 => x"ffffff",
   62281 => x"ffffff",
   62282 => x"ffffff",
   62283 => x"ffffff",
   62284 => x"ffffff",
   62285 => x"ffffff",
   62286 => x"ffffff",
   62287 => x"ffffff",
   62288 => x"ffffff",
   62289 => x"ffffff",
   62290 => x"ffffff",
   62291 => x"ffffff",
   62292 => x"ffffff",
   62293 => x"ffffff",
   62294 => x"ffffff",
   62295 => x"ffffff",
   62296 => x"ffffff",
   62297 => x"ffffff",
   62298 => x"ffffff",
   62299 => x"ffffff",
   62300 => x"ffffff",
   62301 => x"ffffff",
   62302 => x"ffffff",
   62303 => x"ffffff",
   62304 => x"ffffff",
   62305 => x"ffffff",
   62306 => x"ffffff",
   62307 => x"ffffff",
   62308 => x"ffffff",
   62309 => x"ffffff",
   62310 => x"ffffff",
   62311 => x"ffffff",
   62312 => x"ffffff",
   62313 => x"ffffff",
   62314 => x"ffffff",
   62315 => x"ffffff",
   62316 => x"ffffff",
   62317 => x"ffffff",
   62318 => x"ffffff",
   62319 => x"ffffff",
   62320 => x"ffffff",
   62321 => x"ffffff",
   62322 => x"ffffff",
   62323 => x"ffffff",
   62324 => x"ffffff",
   62325 => x"ffffff",
   62326 => x"ffffff",
   62327 => x"ffffff",
   62328 => x"ffffff",
   62329 => x"ffffff",
   62330 => x"ffffff",
   62331 => x"ffffff",
   62332 => x"ffffff",
   62333 => x"ffffff",
   62334 => x"ffffff",
   62335 => x"ffffff",
   62336 => x"ffffff",
   62337 => x"ffffff",
   62338 => x"ffffff",
   62339 => x"ffffff",
   62340 => x"ffffff",
   62341 => x"ffffff",
   62342 => x"ffffff",
   62343 => x"ffffff",
   62344 => x"ffffff",
   62345 => x"ffffff",
   62346 => x"ffffff",
   62347 => x"ffffff",
   62348 => x"ffffff",
   62349 => x"ffffff",
   62350 => x"ffffff",
   62351 => x"ffffff",
   62352 => x"ffffff",
   62353 => x"ffffff",
   62354 => x"ffffff",
   62355 => x"ffffff",
   62356 => x"ffffff",
   62357 => x"ffffff",
   62358 => x"ffffff",
   62359 => x"ffffff",
   62360 => x"ffffff",
   62361 => x"ffffff",
   62362 => x"ffffff",
   62363 => x"ffffff",
   62364 => x"ffffff",
   62365 => x"ffffff",
   62366 => x"ffffff",
   62367 => x"ffffff",
   62368 => x"ffffff",
   62369 => x"ffffff",
   62370 => x"ffffff",
   62371 => x"ffffff",
   62372 => x"ffffff",
   62373 => x"ffffff",
   62374 => x"ffffff",
   62375 => x"ffffff",
   62376 => x"ffffff",
   62377 => x"ffffff",
   62378 => x"ffffff",
   62379 => x"ffffff",
   62380 => x"ffffff",
   62381 => x"ffffff",
   62382 => x"ffffff",
   62383 => x"ffffff",
   62384 => x"ffffff",
   62385 => x"ffffff",
   62386 => x"ffffff",
   62387 => x"ffffff",
   62388 => x"ffffff",
   62389 => x"ffffff",
   62390 => x"ffffff",
   62391 => x"ffffff",
   62392 => x"ffffff",
   62393 => x"ffffff",
   62394 => x"ffffff",
   62395 => x"ffffff",
   62396 => x"ffffff",
   62397 => x"ffffff",
   62398 => x"ffffff",
   62399 => x"ffffff",
   62400 => x"ffffff",
   62401 => x"ffffff",
   62402 => x"ffffff",
   62403 => x"ffffff",
   62404 => x"ffffff",
   62405 => x"ffffff",
   62406 => x"ffffff",
   62407 => x"ffffff",
   62408 => x"ffffff",
   62409 => x"ffffff",
   62410 => x"ffffff",
   62411 => x"ffffff",
   62412 => x"ffffff",
   62413 => x"ffffff",
   62414 => x"ffffff",
   62415 => x"ffffff",
   62416 => x"ffffff",
   62417 => x"ffffff",
   62418 => x"ffffff",
   62419 => x"ffffff",
   62420 => x"ffffff",
   62421 => x"ffffff",
   62422 => x"ffffff",
   62423 => x"ffffff",
   62424 => x"ffffff",
   62425 => x"ffffff",
   62426 => x"ffffff",
   62427 => x"ffffff",
   62428 => x"ffffff",
   62429 => x"ffffff",
   62430 => x"ffffff",
   62431 => x"ffffff",
   62432 => x"ffffff",
   62433 => x"ffffff",
   62434 => x"ffffff",
   62435 => x"ffffff",
   62436 => x"ffffff",
   62437 => x"ffffff",
   62438 => x"ffffff",
   62439 => x"ffffff",
   62440 => x"ffffff",
   62441 => x"ffffff",
   62442 => x"ffffff",
   62443 => x"ffffff",
   62444 => x"ffffff",
   62445 => x"ffffff",
   62446 => x"ffffff",
   62447 => x"ffffff",
   62448 => x"ffffff",
   62449 => x"ffffff",
   62450 => x"ffffff",
   62451 => x"ffffff",
   62452 => x"ffffff",
   62453 => x"ffffff",
   62454 => x"ffffff",
   62455 => x"ffffff",
   62456 => x"ffffff",
   62457 => x"ffffff",
   62458 => x"ffffff",
   62459 => x"ffffff",
   62460 => x"ffffff",
   62461 => x"ffffff",
   62462 => x"ffffff",
   62463 => x"ffffff",
   62464 => x"ffffff",
   62465 => x"ffffff",
   62466 => x"ffffff",
   62467 => x"ffffff",
   62468 => x"ffffff",
   62469 => x"ffffff",
   62470 => x"ffffff",
   62471 => x"ffffff",
   62472 => x"ffffff",
   62473 => x"ffffff",
   62474 => x"ffffff",
   62475 => x"ffffff",
   62476 => x"ffffff",
   62477 => x"ffffff",
   62478 => x"ffffff",
   62479 => x"ffffff",
   62480 => x"ffffff",
   62481 => x"ffffff",
   62482 => x"ffffff",
   62483 => x"ffffff",
   62484 => x"ffffff",
   62485 => x"ffffff",
   62486 => x"ffffff",
   62487 => x"ffffff",
   62488 => x"ffffff",
   62489 => x"ffffff",
   62490 => x"ffffff",
   62491 => x"ffffff",
   62492 => x"ffffff",
   62493 => x"ffffff",
   62494 => x"ffffff",
   62495 => x"ffffff",
   62496 => x"ffffff",
   62497 => x"ffffff",
   62498 => x"ffffff",
   62499 => x"ffffff",
   62500 => x"ffffff",
   62501 => x"ffffff",
   62502 => x"ffffff",
   62503 => x"ffffff",
   62504 => x"ffffff",
   62505 => x"ffffff",
   62506 => x"ffffff",
   62507 => x"ffffff",
   62508 => x"ffffff",
   62509 => x"ffffff",
   62510 => x"ffffff",
   62511 => x"ffffff",
   62512 => x"ffffff",
   62513 => x"ffffff",
   62514 => x"ffffff",
   62515 => x"ffffff",
   62516 => x"ffffff",
   62517 => x"ffffff",
   62518 => x"ffffff",
   62519 => x"ffffff",
   62520 => x"ffffff",
   62521 => x"ffffff",
   62522 => x"ffffff",
   62523 => x"ffffff",
   62524 => x"ffffff",
   62525 => x"ffffff",
   62526 => x"ffffff",
   62527 => x"ffffff",
   62528 => x"ffffff",
   62529 => x"ffffff",
   62530 => x"ffffff",
   62531 => x"ffffff",
   62532 => x"ffffff",
   62533 => x"ffffff",
   62534 => x"ffffff",
   62535 => x"ffffff",
   62536 => x"ffffff",
   62537 => x"ffffff",
   62538 => x"ffffff",
   62539 => x"ffffff",
   62540 => x"ffffff",
   62541 => x"ffffff",
   62542 => x"ffffff",
   62543 => x"ffffff",
   62544 => x"ffffff",
   62545 => x"ffffff",
   62546 => x"ffffff",
   62547 => x"ffffff",
   62548 => x"ffffff",
   62549 => x"ffffff",
   62550 => x"ffffff",
   62551 => x"ffffff",
   62552 => x"ffffff",
   62553 => x"ffffff",
   62554 => x"ffffff",
   62555 => x"ffffff",
   62556 => x"ffffff",
   62557 => x"ffffff",
   62558 => x"ffffff",
   62559 => x"ffffff",
   62560 => x"ffffff",
   62561 => x"ffffff",
   62562 => x"ffffff",
   62563 => x"ffffff",
   62564 => x"ffffff",
   62565 => x"ffffff",
   62566 => x"ffffff",
   62567 => x"ffffff",
   62568 => x"ffffff",
   62569 => x"ffffff",
   62570 => x"ffffff",
   62571 => x"ffffff",
   62572 => x"ffffff",
   62573 => x"ffffff",
   62574 => x"ffffff",
   62575 => x"ffffff",
   62576 => x"ffffff",
   62577 => x"ffffff",
   62578 => x"ffffff",
   62579 => x"ffffff",
   62580 => x"ffffff",
   62581 => x"ffffff",
   62582 => x"ffffff",
   62583 => x"ffffff",
   62584 => x"ffffff",
   62585 => x"ffffff",
   62586 => x"ffffff",
   62587 => x"ffffff",
   62588 => x"ffffff",
   62589 => x"ffffff",
   62590 => x"ffffff",
   62591 => x"ffffff",
   62592 => x"ffffff",
   62593 => x"ffffff",
   62594 => x"ffffff",
   62595 => x"ffffff",
   62596 => x"ffffff",
   62597 => x"ffffff",
   62598 => x"ffffff",
   62599 => x"ffffff",
   62600 => x"ffffff",
   62601 => x"ffffff",
   62602 => x"ffffff",
   62603 => x"ffffff",
   62604 => x"ffffff",
   62605 => x"ffffff",
   62606 => x"ffffff",
   62607 => x"ffffff",
   62608 => x"ffffff",
   62609 => x"ffffff",
   62610 => x"ffffff",
   62611 => x"ffffff",
   62612 => x"ffffff",
   62613 => x"ffffff",
   62614 => x"ffffff",
   62615 => x"ffffff",
   62616 => x"ffffff",
   62617 => x"ffffff",
   62618 => x"ffffff",
   62619 => x"ffffff",
   62620 => x"ffffff",
   62621 => x"ffffff",
   62622 => x"ffffff",
   62623 => x"ffffff",
   62624 => x"ffffff",
   62625 => x"ffffff",
   62626 => x"ffffff",
   62627 => x"ffffff",
   62628 => x"ffffff",
   62629 => x"ffffff",
   62630 => x"ffffff",
   62631 => x"ffffff",
   62632 => x"ffffff",
   62633 => x"ffffff",
   62634 => x"ffffff",
   62635 => x"ffffff",
   62636 => x"ffffff",
   62637 => x"ffffff",
   62638 => x"ffffff",
   62639 => x"ffffff",
   62640 => x"ffffff",
   62641 => x"ffffff",
   62642 => x"ffffff",
   62643 => x"ffffff",
   62644 => x"ffffff",
   62645 => x"ffffff",
   62646 => x"ffffff",
   62647 => x"ffffff",
   62648 => x"ffffff",
   62649 => x"ffffff",
   62650 => x"ffffff",
   62651 => x"ffffff",
   62652 => x"ffffff",
   62653 => x"ffffff",
   62654 => x"ffffff",
   62655 => x"ffffff",
   62656 => x"ffffff",
   62657 => x"ffffff",
   62658 => x"ffffff",
   62659 => x"ffffff",
   62660 => x"ffffff",
   62661 => x"ffffff",
   62662 => x"ffffff",
   62663 => x"ffffff",
   62664 => x"ffffff",
   62665 => x"ffffff",
   62666 => x"ffffff",
   62667 => x"ffffff",
   62668 => x"ffffff",
   62669 => x"ffffff",
   62670 => x"ffffff",
   62671 => x"ffffff",
   62672 => x"ffffff",
   62673 => x"ffffff",
   62674 => x"ffffff",
   62675 => x"ffffff",
   62676 => x"ffffff",
   62677 => x"ffffff",
   62678 => x"ffffff",
   62679 => x"ffffff",
   62680 => x"ffffff",
   62681 => x"ffffff",
   62682 => x"ffffff",
   62683 => x"ffffff",
   62684 => x"ffffff",
   62685 => x"ffffff",
   62686 => x"ffffff",
   62687 => x"ffffff",
   62688 => x"ffffff",
   62689 => x"ffffff",
   62690 => x"ffffff",
   62691 => x"ffffff",
   62692 => x"ffffff",
   62693 => x"ffffff",
   62694 => x"ffffff",
   62695 => x"ffffff",
   62696 => x"ffffff",
   62697 => x"ffffff",
   62698 => x"ffffff",
   62699 => x"ffffff",
   62700 => x"ffffff",
   62701 => x"ffffff",
   62702 => x"ffffff",
   62703 => x"ffffff",
   62704 => x"ffffff",
   62705 => x"ffffff",
   62706 => x"ffffff",
   62707 => x"ffffff",
   62708 => x"ffffff",
   62709 => x"ffffff",
   62710 => x"ffffff",
   62711 => x"ffffff",
   62712 => x"ffffff",
   62713 => x"ffffff",
   62714 => x"ffffff",
   62715 => x"ffffff",
   62716 => x"ffffff",
   62717 => x"ffffff",
   62718 => x"ffffff",
   62719 => x"ffffff",
   62720 => x"ffffff",
   62721 => x"ffffff",
   62722 => x"ffffff",
   62723 => x"ffffff",
   62724 => x"ffffff",
   62725 => x"ffffff",
   62726 => x"ffffff",
   62727 => x"ffffff",
   62728 => x"ffffff",
   62729 => x"ffffff",
   62730 => x"ffffff",
   62731 => x"ffffff",
   62732 => x"ffffff",
   62733 => x"ffffff",
   62734 => x"ffffff",
   62735 => x"ffffff",
   62736 => x"ffffff",
   62737 => x"ffffff",
   62738 => x"ffffff",
   62739 => x"ffffff",
   62740 => x"ffffff",
   62741 => x"ffffff",
   62742 => x"ffffff",
   62743 => x"ffffff",
   62744 => x"ffffff",
   62745 => x"ffffff",
   62746 => x"ffffff",
   62747 => x"ffffff",
   62748 => x"ffffff",
   62749 => x"ffffff",
   62750 => x"ffffff",
   62751 => x"ffffff",
   62752 => x"ffffff",
   62753 => x"ffffff",
   62754 => x"ffffff",
   62755 => x"ffffff",
   62756 => x"ffffff",
   62757 => x"ffffff",
   62758 => x"ffffff",
   62759 => x"ffffff",
   62760 => x"ffffff",
   62761 => x"ffffff",
   62762 => x"ffffff",
   62763 => x"ffffff",
   62764 => x"ffffff",
   62765 => x"ffffff",
   62766 => x"ffffff",
   62767 => x"ffffff",
   62768 => x"ffffff",
   62769 => x"ffffff",
   62770 => x"ffffff",
   62771 => x"ffffff",
   62772 => x"ffffff",
   62773 => x"ffffff",
   62774 => x"ffffff",
   62775 => x"ffffff",
   62776 => x"ffffff",
   62777 => x"ffffff",
   62778 => x"ffffff",
   62779 => x"ffffff",
   62780 => x"ffffff",
   62781 => x"ffffff",
   62782 => x"ffffff",
   62783 => x"ffffff",
   62784 => x"ffffff",
   62785 => x"ffffff",
   62786 => x"ffffff",
   62787 => x"ffffff",
   62788 => x"ffffff",
   62789 => x"ffffff",
   62790 => x"ffffff",
   62791 => x"ffffff",
   62792 => x"ffffff",
   62793 => x"ffffff",
   62794 => x"ffffff",
   62795 => x"ffffff",
   62796 => x"ffffff",
   62797 => x"ffffff",
   62798 => x"ffffff",
   62799 => x"ffffff",
   62800 => x"ffffff",
   62801 => x"ffffff",
   62802 => x"ffffff",
   62803 => x"ffffff",
   62804 => x"ffffff",
   62805 => x"ffffff",
   62806 => x"ffffff",
   62807 => x"ffffff",
   62808 => x"ffffff",
   62809 => x"ffffff",
   62810 => x"ffffff",
   62811 => x"ffffff",
   62812 => x"ffffff",
   62813 => x"ffffff",
   62814 => x"ffffff",
   62815 => x"ffffff",
   62816 => x"ffffff",
   62817 => x"ffffff",
   62818 => x"ffffff",
   62819 => x"ffffff",
   62820 => x"ffffff",
   62821 => x"ffffff",
   62822 => x"ffffff",
   62823 => x"ffffff",
   62824 => x"ffffff",
   62825 => x"ffffff",
   62826 => x"ffffff",
   62827 => x"ffffff",
   62828 => x"ffffff",
   62829 => x"ffffff",
   62830 => x"ffffff",
   62831 => x"ffffff",
   62832 => x"ffffff",
   62833 => x"ffffff",
   62834 => x"ffffff",
   62835 => x"ffffff",
   62836 => x"ffffff",
   62837 => x"ffffff",
   62838 => x"ffffff",
   62839 => x"ffffff",
   62840 => x"ffffff",
   62841 => x"ffffff",
   62842 => x"ffffff",
   62843 => x"ffffff",
   62844 => x"ffffff",
   62845 => x"ffffff",
   62846 => x"ffffff",
   62847 => x"ffffff",
   62848 => x"ffffff",
   62849 => x"ffffff",
   62850 => x"ffffff",
   62851 => x"ffffff",
   62852 => x"ffffff",
   62853 => x"ffffff",
   62854 => x"ffffff",
   62855 => x"ffffff",
   62856 => x"ffffff",
   62857 => x"ffffff",
   62858 => x"ffffff",
   62859 => x"ffffff",
   62860 => x"ffffff",
   62861 => x"ffffff",
   62862 => x"ffffff",
   62863 => x"ffffff",
   62864 => x"ffffff",
   62865 => x"ffffff",
   62866 => x"ffffff",
   62867 => x"ffffff",
   62868 => x"ffffff",
   62869 => x"ffffff",
   62870 => x"ffffff",
   62871 => x"ffffff",
   62872 => x"ffffff",
   62873 => x"ffffff",
   62874 => x"ffffff",
   62875 => x"ffffff",
   62876 => x"ffffff",
   62877 => x"ffffff",
   62878 => x"ffffff",
   62879 => x"ffffff",
   62880 => x"ffffff",
   62881 => x"ffffff",
   62882 => x"ffffff",
   62883 => x"ffffff",
   62884 => x"ffffff",
   62885 => x"ffffff",
   62886 => x"ffffff",
   62887 => x"ffffff",
   62888 => x"ffffff",
   62889 => x"ffffff",
   62890 => x"ffffff",
   62891 => x"ffffff",
   62892 => x"ffffff",
   62893 => x"ffffff",
   62894 => x"ffffff",
   62895 => x"ffffff",
   62896 => x"ffffff",
   62897 => x"ffffff",
   62898 => x"ffffff",
   62899 => x"ffffff",
   62900 => x"ffffff",
   62901 => x"ffffff",
   62902 => x"ffffff",
   62903 => x"ffffff",
   62904 => x"ffffff",
   62905 => x"ffffff",
   62906 => x"ffffff",
   62907 => x"ffffff",
   62908 => x"ffffff",
   62909 => x"ffffff",
   62910 => x"ffffff",
   62911 => x"ffffff",
   62912 => x"ffffff",
   62913 => x"ffffff",
   62914 => x"ffffff",
   62915 => x"ffffff",
   62916 => x"ffffff",
   62917 => x"ffffff",
   62918 => x"ffffff",
   62919 => x"ffffff",
   62920 => x"ffffff",
   62921 => x"ffffff",
   62922 => x"ffffff",
   62923 => x"ffffff",
   62924 => x"ffffff",
   62925 => x"ffffff",
   62926 => x"ffffff",
   62927 => x"ffffff",
   62928 => x"ffffff",
   62929 => x"ffffff",
   62930 => x"ffffff",
   62931 => x"ffffff",
   62932 => x"ffffff",
   62933 => x"ffffff",
   62934 => x"ffffff",
   62935 => x"ffffff",
   62936 => x"ffffff",
   62937 => x"ffffff",
   62938 => x"ffffff",
   62939 => x"ffffff",
   62940 => x"ffffff",
   62941 => x"ffffff",
   62942 => x"ffffff",
   62943 => x"ffffff",
   62944 => x"ffffff",
   62945 => x"ffffff",
   62946 => x"ffffff",
   62947 => x"ffffff",
   62948 => x"ffffff",
   62949 => x"ffffff",
   62950 => x"ffffff",
   62951 => x"ffffff",
   62952 => x"ffffff",
   62953 => x"ffffff",
   62954 => x"ffffff",
   62955 => x"ffffff",
   62956 => x"ffffff",
   62957 => x"ffffff",
   62958 => x"ffffff",
   62959 => x"ffffff",
   62960 => x"ffffff",
   62961 => x"ffffff",
   62962 => x"ffffff",
   62963 => x"ffffff",
   62964 => x"ffffff",
   62965 => x"ffffff",
   62966 => x"ffffff",
   62967 => x"ffffff",
   62968 => x"ffffff",
   62969 => x"ffffff",
   62970 => x"ffffff",
   62971 => x"ffffff",
   62972 => x"ffffff",
   62973 => x"ffffff",
   62974 => x"ffffff",
   62975 => x"ffffff",
   62976 => x"ffffff",
   62977 => x"ffffff",
   62978 => x"ffffff",
   62979 => x"ffffff",
   62980 => x"ffffff",
   62981 => x"ffffff",
   62982 => x"ffffff",
   62983 => x"ffffff",
   62984 => x"ffffff",
   62985 => x"ffffff",
   62986 => x"ffffff",
   62987 => x"ffffff",
   62988 => x"ffffff",
   62989 => x"ffffff",
   62990 => x"ffffff",
   62991 => x"ffffff",
   62992 => x"ffffff",
   62993 => x"ffffff",
   62994 => x"ffffff",
   62995 => x"ffffff",
   62996 => x"ffffff",
   62997 => x"ffffff",
   62998 => x"ffffff",
   62999 => x"ffffff",
   63000 => x"ffffff",
   63001 => x"ffffff",
   63002 => x"ffffff",
   63003 => x"ffffff",
   63004 => x"ffffff",
   63005 => x"ffffff",
   63006 => x"ffffff",
   63007 => x"ffffff",
   63008 => x"ffffff",
   63009 => x"ffffff",
   63010 => x"ffffff",
   63011 => x"ffffff",
   63012 => x"ffffff",
   63013 => x"ffffff",
   63014 => x"ffffff",
   63015 => x"ffffff",
   63016 => x"ffffff",
   63017 => x"ffffff",
   63018 => x"ffffff",
   63019 => x"ffffff",
   63020 => x"ffffff",
   63021 => x"ffffff",
   63022 => x"ffffff",
   63023 => x"ffffff",
   63024 => x"ffffff",
   63025 => x"ffffff",
   63026 => x"ffffff",
   63027 => x"ffffff",
   63028 => x"ffffff",
   63029 => x"ffffff",
   63030 => x"ffffff",
   63031 => x"ffffff",
   63032 => x"ffffff",
   63033 => x"ffffff",
   63034 => x"ffffff",
   63035 => x"ffffff",
   63036 => x"ffffff",
   63037 => x"ffffff",
   63038 => x"ffffff",
   63039 => x"ffffff",
   63040 => x"ffffff",
   63041 => x"ffffff",
   63042 => x"ffffff",
   63043 => x"ffffff",
   63044 => x"ffffff",
   63045 => x"ffffff",
   63046 => x"ffffff",
   63047 => x"ffffff",
   63048 => x"ffffff",
   63049 => x"ffffff",
   63050 => x"ffffff",
   63051 => x"ffffff",
   63052 => x"ffffff",
   63053 => x"ffffff",
   63054 => x"ffffff",
   63055 => x"ffffff",
   63056 => x"ffffff",
   63057 => x"ffffff",
   63058 => x"ffffff",
   63059 => x"ffffff",
   63060 => x"ffffff",
   63061 => x"ffffff",
   63062 => x"ffffff",
   63063 => x"ffffff",
   63064 => x"ffffff",
   63065 => x"ffffff",
   63066 => x"ffffff",
   63067 => x"ffffff",
   63068 => x"ffffff",
   63069 => x"ffffff",
   63070 => x"ffffff",
   63071 => x"ffffff",
   63072 => x"ffffff",
   63073 => x"ffffff",
   63074 => x"ffffff",
   63075 => x"ffffff",
   63076 => x"ffffff",
   63077 => x"ffffff",
   63078 => x"ffffff",
   63079 => x"ffffff",
   63080 => x"ffffff",
   63081 => x"ffffff",
   63082 => x"ffffff",
   63083 => x"ffffff",
   63084 => x"ffffff",
   63085 => x"ffffff",
   63086 => x"ffffff",
   63087 => x"ffffff",
   63088 => x"ffffff",
   63089 => x"ffffff",
   63090 => x"ffffff",
   63091 => x"ffffff",
   63092 => x"ffffff",
   63093 => x"ffffff",
   63094 => x"ffffff",
   63095 => x"ffffff",
   63096 => x"ffffff",
   63097 => x"ffffff",
   63098 => x"ffffff",
   63099 => x"ffffff",
   63100 => x"ffffff",
   63101 => x"ffffff",
   63102 => x"ffffff",
   63103 => x"ffffff",
   63104 => x"ffffff",
   63105 => x"ffffff",
   63106 => x"ffffff",
   63107 => x"ffffff",
   63108 => x"ffffff",
   63109 => x"ffffff",
   63110 => x"ffffff",
   63111 => x"ffffff",
   63112 => x"ffffff",
   63113 => x"ffffff",
   63114 => x"ffffff",
   63115 => x"ffffff",
   63116 => x"ffffff",
   63117 => x"ffffff",
   63118 => x"ffffff",
   63119 => x"ffffff",
   63120 => x"ffffff",
   63121 => x"ffffff",
   63122 => x"ffffff",
   63123 => x"ffffff",
   63124 => x"ffffff",
   63125 => x"ffffff",
   63126 => x"ffffff",
   63127 => x"ffffff",
   63128 => x"ffffff",
   63129 => x"ffffff",
   63130 => x"ffffff",
   63131 => x"ffffff",
   63132 => x"ffffff",
   63133 => x"ffffff",
   63134 => x"ffffff",
   63135 => x"ffffff",
   63136 => x"ffffff",
   63137 => x"ffffff",
   63138 => x"ffffff",
   63139 => x"ffffff",
   63140 => x"ffffff",
   63141 => x"ffffff",
   63142 => x"ffffff",
   63143 => x"ffffff",
   63144 => x"ffffff",
   63145 => x"ffffff",
   63146 => x"ffffff",
   63147 => x"ffffff",
   63148 => x"ffffff",
   63149 => x"ffffff",
   63150 => x"ffffff",
   63151 => x"ffffff",
   63152 => x"ffffff",
   63153 => x"ffffff",
   63154 => x"ffffff",
   63155 => x"ffffff",
   63156 => x"ffffff",
   63157 => x"ffffff",
   63158 => x"ffffff",
   63159 => x"ffffff",
   63160 => x"ffffff",
   63161 => x"ffffff",
   63162 => x"ffffff",
   63163 => x"ffffff",
   63164 => x"ffffff",
   63165 => x"ffffff",
   63166 => x"ffffff",
   63167 => x"ffffff",
   63168 => x"ffffff",
   63169 => x"ffffff",
   63170 => x"ffffff",
   63171 => x"ffffff",
   63172 => x"ffffff",
   63173 => x"ffffff",
   63174 => x"ffffff",
   63175 => x"ffffff",
   63176 => x"ffffff",
   63177 => x"ffffff",
   63178 => x"ffffff",
   63179 => x"ffffff",
   63180 => x"ffffff",
   63181 => x"ffffff",
   63182 => x"ffffff",
   63183 => x"ffffff",
   63184 => x"ffffff",
   63185 => x"ffffff",
   63186 => x"ffffff",
   63187 => x"ffffff",
   63188 => x"ffffff",
   63189 => x"ffffff",
   63190 => x"ffffff",
   63191 => x"ffffff",
   63192 => x"ffffff",
   63193 => x"ffffff",
   63194 => x"ffffff",
   63195 => x"ffffff",
   63196 => x"ffffff",
   63197 => x"ffffff",
   63198 => x"ffffff",
   63199 => x"ffffff",
   63200 => x"ffffff",
   63201 => x"ffffff",
   63202 => x"ffffff",
   63203 => x"ffffff",
   63204 => x"ffffff",
   63205 => x"ffffff",
   63206 => x"ffffff",
   63207 => x"ffffff",
   63208 => x"ffffff",
   63209 => x"ffffff",
   63210 => x"ffffff",
   63211 => x"ffffff",
   63212 => x"ffffff",
   63213 => x"ffffff",
   63214 => x"ffffff",
   63215 => x"ffffff",
   63216 => x"ffffff",
   63217 => x"ffffff",
   63218 => x"ffffff",
   63219 => x"ffffff",
   63220 => x"ffffff",
   63221 => x"ffffff",
   63222 => x"ffffff",
   63223 => x"ffffff",
   63224 => x"ffffff",
   63225 => x"ffffff",
   63226 => x"ffffff",
   63227 => x"ffffff",
   63228 => x"ffffff",
   63229 => x"ffffff",
   63230 => x"ffffff",
   63231 => x"ffffff",
   63232 => x"ffffff",
   63233 => x"ffffff",
   63234 => x"ffffff",
   63235 => x"ffffff",
   63236 => x"ffffff",
   63237 => x"ffffff",
   63238 => x"ffffff",
   63239 => x"ffffff",
   63240 => x"ffffff",
   63241 => x"ffffff",
   63242 => x"ffffff",
   63243 => x"ffffff",
   63244 => x"ffffff",
   63245 => x"ffffff",
   63246 => x"ffffff",
   63247 => x"ffffff",
   63248 => x"ffffff",
   63249 => x"ffffff",
   63250 => x"ffffff",
   63251 => x"ffffff",
   63252 => x"ffffff",
   63253 => x"ffffff",
   63254 => x"ffffff",
   63255 => x"ffffff",
   63256 => x"ffffff",
   63257 => x"ffffff",
   63258 => x"ffffff",
   63259 => x"ffffff",
   63260 => x"ffffff",
   63261 => x"ffffff",
   63262 => x"ffffff",
   63263 => x"ffffff",
   63264 => x"ffffff",
   63265 => x"ffffff",
   63266 => x"ffffff",
   63267 => x"ffffff",
   63268 => x"ffffff",
   63269 => x"ffffff",
   63270 => x"ffffff",
   63271 => x"ffffff",
   63272 => x"ffffff",
   63273 => x"ffffff",
   63274 => x"ffffff",
   63275 => x"ffffff",
   63276 => x"ffffff",
   63277 => x"ffffff",
   63278 => x"ffffff",
   63279 => x"ffffff",
   63280 => x"ffffff",
   63281 => x"ffffff",
   63282 => x"ffffff",
   63283 => x"ffffff",
   63284 => x"ffffff",
   63285 => x"ffffff",
   63286 => x"ffffff",
   63287 => x"ffffff",
   63288 => x"ffffff",
   63289 => x"ffffff",
   63290 => x"ffffff",
   63291 => x"ffffff",
   63292 => x"ffffff",
   63293 => x"ffffff",
   63294 => x"ffffff",
   63295 => x"ffffff",
   63296 => x"ffffff",
   63297 => x"ffffff",
   63298 => x"ffffff",
   63299 => x"ffffff",
   63300 => x"ffffff",
   63301 => x"ffffff",
   63302 => x"ffffff",
   63303 => x"ffffff",
   63304 => x"ffffff",
   63305 => x"ffffff",
   63306 => x"ffffff",
   63307 => x"ffffff",
   63308 => x"ffffff",
   63309 => x"ffffff",
   63310 => x"ffffff",
   63311 => x"ffffff",
   63312 => x"ffffff",
   63313 => x"ffffff",
   63314 => x"ffffff",
   63315 => x"ffffff",
   63316 => x"ffffff",
   63317 => x"ffffff",
   63318 => x"ffffff",
   63319 => x"ffffff",
   63320 => x"ffffff",
   63321 => x"ffffff",
   63322 => x"ffffff",
   63323 => x"ffffff",
   63324 => x"ffffff",
   63325 => x"ffffff",
   63326 => x"ffffff",
   63327 => x"ffffff",
   63328 => x"ffffff",
   63329 => x"ffffff",
   63330 => x"ffffff",
   63331 => x"ffffff",
   63332 => x"ffffff",
   63333 => x"ffffff",
   63334 => x"ffffff",
   63335 => x"ffffff",
   63336 => x"ffffff",
   63337 => x"ffffff",
   63338 => x"ffffff",
   63339 => x"ffffff",
   63340 => x"ffffff",
   63341 => x"ffffff",
   63342 => x"ffffff",
   63343 => x"ffffff",
   63344 => x"ffffff",
   63345 => x"ffffff",
   63346 => x"ffffff",
   63347 => x"ffffff",
   63348 => x"ffffff",
   63349 => x"ffffff",
   63350 => x"ffffff",
   63351 => x"ffffff",
   63352 => x"ffffff",
   63353 => x"ffffff",
   63354 => x"ffffff",
   63355 => x"ffffff",
   63356 => x"ffffff",
   63357 => x"ffffff",
   63358 => x"ffffff",
   63359 => x"ffffff",
   63360 => x"ffffff",
   63361 => x"ffffff",
   63362 => x"ffffff",
   63363 => x"ffffff",
   63364 => x"ffffff",
   63365 => x"ffffff",
   63366 => x"ffffff",
   63367 => x"ffffff",
   63368 => x"ffffff",
   63369 => x"ffffff",
   63370 => x"ffffff",
   63371 => x"ffffff",
   63372 => x"ffffff",
   63373 => x"ffffff",
   63374 => x"ffffff",
   63375 => x"ffffff",
   63376 => x"ffffff",
   63377 => x"ffffff",
   63378 => x"ffffff",
   63379 => x"ffffff",
   63380 => x"ffffff",
   63381 => x"ffffff",
   63382 => x"ffffff",
   63383 => x"ffffff",
   63384 => x"ffffff",
   63385 => x"ffffff",
   63386 => x"ffffff",
   63387 => x"ffffff",
   63388 => x"ffffff",
   63389 => x"ffffff",
   63390 => x"ffffff",
   63391 => x"ffffff",
   63392 => x"ffffff",
   63393 => x"ffffff",
   63394 => x"ffffff",
   63395 => x"ffffff",
   63396 => x"ffffff",
   63397 => x"ffffff",
   63398 => x"ffffff",
   63399 => x"ffffff",
   63400 => x"ffffff",
   63401 => x"ffffff",
   63402 => x"ffffff",
   63403 => x"ffffff",
   63404 => x"ffffff",
   63405 => x"ffffff",
   63406 => x"ffffff",
   63407 => x"ffffff",
   63408 => x"ffffff",
   63409 => x"ffffff",
   63410 => x"ffffff",
   63411 => x"ffffff",
   63412 => x"ffffff",
   63413 => x"ffffff",
   63414 => x"ffffff",
   63415 => x"ffffff",
   63416 => x"ffffff",
   63417 => x"ffffff",
   63418 => x"ffffff",
   63419 => x"ffffff",
   63420 => x"ffffff",
   63421 => x"ffffff",
   63422 => x"ffffff",
   63423 => x"ffffff",
   63424 => x"ffffff",
   63425 => x"ffffff",
   63426 => x"ffffff",
   63427 => x"ffffff",
   63428 => x"ffffff",
   63429 => x"ffffff",
   63430 => x"ffffff",
   63431 => x"ffffff",
   63432 => x"ffffff",
   63433 => x"ffffff",
   63434 => x"ffffff",
   63435 => x"ffffff",
   63436 => x"ffffff",
   63437 => x"ffffff",
   63438 => x"ffffff",
   63439 => x"ffffff",
   63440 => x"ffffff",
   63441 => x"ffffff",
   63442 => x"ffffff",
   63443 => x"ffffff",
   63444 => x"ffffff",
   63445 => x"ffffff",
   63446 => x"ffffff",
   63447 => x"ffffff",
   63448 => x"ffffff",
   63449 => x"ffffff",
   63450 => x"ffffff",
   63451 => x"ffffff",
   63452 => x"ffffff",
   63453 => x"ffffff",
   63454 => x"ffffff",
   63455 => x"ffffff",
   63456 => x"ffffff",
   63457 => x"ffffff",
   63458 => x"ffffff",
   63459 => x"ffffff",
   63460 => x"ffffff",
   63461 => x"ffffff",
   63462 => x"ffffff",
   63463 => x"ffffff",
   63464 => x"ffffff",
   63465 => x"ffffff",
   63466 => x"ffffff",
   63467 => x"ffffff",
   63468 => x"ffffff",
   63469 => x"ffffff",
   63470 => x"ffffff",
   63471 => x"ffffff",
   63472 => x"ffffff",
   63473 => x"ffffff",
   63474 => x"ffffff",
   63475 => x"ffffff",
   63476 => x"ffffff",
   63477 => x"ffffff",
   63478 => x"ffffff",
   63479 => x"ffffff",
   63480 => x"ffffff",
   63481 => x"ffffff",
   63482 => x"ffffff",
   63483 => x"ffffff",
   63484 => x"ffffff",
   63485 => x"ffffff",
   63486 => x"ffffff",
   63487 => x"ffffff",
   63488 => x"ffffff",
   63489 => x"ffffff",
   63490 => x"ffffff",
   63491 => x"ffffff",
   63492 => x"ffffff",
   63493 => x"ffffff",
   63494 => x"ffffff",
   63495 => x"ffffff",
   63496 => x"ffffff",
   63497 => x"ffffff",
   63498 => x"ffffff",
   63499 => x"ffffff",
   63500 => x"ffffff",
   63501 => x"ffffff",
   63502 => x"ffffff",
   63503 => x"ffffff",
   63504 => x"ffffff",
   63505 => x"ffffff",
   63506 => x"ffffff",
   63507 => x"ffffff",
   63508 => x"ffffff",
   63509 => x"ffffff",
   63510 => x"ffffff",
   63511 => x"ffffff",
   63512 => x"ffffff",
   63513 => x"ffffff",
   63514 => x"ffffff",
   63515 => x"ffffff",
   63516 => x"ffffff",
   63517 => x"ffffff",
   63518 => x"ffffff",
   63519 => x"ffffff",
   63520 => x"ffffff",
   63521 => x"ffffff",
   63522 => x"ffffff",
   63523 => x"ffffff",
   63524 => x"ffffff",
   63525 => x"ffffff",
   63526 => x"ffffff",
   63527 => x"ffffff",
   63528 => x"ffffff",
   63529 => x"ffffff",
   63530 => x"ffffff",
   63531 => x"ffffff",
   63532 => x"ffffff",
   63533 => x"ffffff",
   63534 => x"ffffff",
   63535 => x"ffffff",
   63536 => x"ffffff",
   63537 => x"ffffff",
   63538 => x"ffffff",
   63539 => x"ffffff",
   63540 => x"ffffff",
   63541 => x"ffffff",
   63542 => x"ffffff",
   63543 => x"ffffff",
   63544 => x"ffffff",
   63545 => x"ffffff",
   63546 => x"ffffff",
   63547 => x"ffffff",
   63548 => x"ffffff",
   63549 => x"ffffff",
   63550 => x"ffffff",
   63551 => x"ffffff",
   63552 => x"ffffff",
   63553 => x"ffffff",
   63554 => x"ffffff",
   63555 => x"ffffff",
   63556 => x"ffffff",
   63557 => x"ffffff",
   63558 => x"ffffff",
   63559 => x"ffffff",
   63560 => x"ffffff",
   63561 => x"ffffff",
   63562 => x"ffffff",
   63563 => x"ffffff",
   63564 => x"ffffff",
   63565 => x"ffffff",
   63566 => x"ffffff",
   63567 => x"ffffff",
   63568 => x"ffffff",
   63569 => x"ffffff",
   63570 => x"ffffff",
   63571 => x"ffffff",
   63572 => x"ffffff",
   63573 => x"ffffff",
   63574 => x"ffffff",
   63575 => x"ffffff",
   63576 => x"ffffff",
   63577 => x"ffffff",
   63578 => x"ffffff",
   63579 => x"ffffff",
   63580 => x"ffffff",
   63581 => x"ffffff",
   63582 => x"ffffff",
   63583 => x"ffffff",
   63584 => x"ffffff",
   63585 => x"ffffff",
   63586 => x"ffffff",
   63587 => x"ffffff",
   63588 => x"ffffff",
   63589 => x"ffffff",
   63590 => x"ffffff",
   63591 => x"ffffff",
   63592 => x"ffffff",
   63593 => x"ffffff",
   63594 => x"ffffff",
   63595 => x"ffffff",
   63596 => x"ffffff",
   63597 => x"ffffff",
   63598 => x"ffffff",
   63599 => x"ffffff",
   63600 => x"ffffff",
   63601 => x"ffffff",
   63602 => x"ffffff",
   63603 => x"ffffff",
   63604 => x"ffffff",
   63605 => x"ffffff",
   63606 => x"ffffff",
   63607 => x"ffffff",
   63608 => x"ffffff",
   63609 => x"ffffff",
   63610 => x"ffffff",
   63611 => x"ffffff",
   63612 => x"ffffff",
   63613 => x"ffffff",
   63614 => x"ffffff",
   63615 => x"ffffff",
   63616 => x"ffffff",
   63617 => x"ffffff",
   63618 => x"ffffff",
   63619 => x"ffffff",
   63620 => x"ffffff",
   63621 => x"ffffff",
   63622 => x"ffffff",
   63623 => x"ffffff",
   63624 => x"ffffff",
   63625 => x"ffffff",
   63626 => x"ffffff",
   63627 => x"ffffff",
   63628 => x"ffffff",
   63629 => x"ffffff",
   63630 => x"ffffff",
   63631 => x"ffffff",
   63632 => x"ffffff",
   63633 => x"ffffff",
   63634 => x"ffffff",
   63635 => x"ffffff",
   63636 => x"ffffff",
   63637 => x"ffffff",
   63638 => x"ffffff",
   63639 => x"ffffff",
   63640 => x"ffffff",
   63641 => x"ffffff",
   63642 => x"ffffff",
   63643 => x"ffffff",
   63644 => x"ffffff",
   63645 => x"ffffff",
   63646 => x"ffffff",
   63647 => x"ffffff",
   63648 => x"ffffff",
   63649 => x"ffffff",
   63650 => x"ffffff",
   63651 => x"ffffff",
   63652 => x"ffffff",
   63653 => x"ffffff",
   63654 => x"ffffff",
   63655 => x"ffffff",
   63656 => x"ffffff",
   63657 => x"ffffff",
   63658 => x"ffffff",
   63659 => x"ffffff",
   63660 => x"ffffff",
   63661 => x"ffffff",
   63662 => x"ffffff",
   63663 => x"ffffff",
   63664 => x"ffffff",
   63665 => x"ffffff",
   63666 => x"ffffff",
   63667 => x"ffffff",
   63668 => x"ffffff",
   63669 => x"ffffff",
   63670 => x"ffffff",
   63671 => x"ffffff",
   63672 => x"ffffff",
   63673 => x"ffffff",
   63674 => x"ffffff",
   63675 => x"ffffff",
   63676 => x"ffffff",
   63677 => x"ffffff",
   63678 => x"ffffff",
   63679 => x"ffffff",
   63680 => x"ffffff",
   63681 => x"ffffff",
   63682 => x"ffffff",
   63683 => x"ffffff",
   63684 => x"ffffff",
   63685 => x"ffffff",
   63686 => x"ffffff",
   63687 => x"ffffff",
   63688 => x"ffffff",
   63689 => x"ffffff",
   63690 => x"ffffff",
   63691 => x"ffffff",
   63692 => x"ffffff",
   63693 => x"ffffff",
   63694 => x"ffffff",
   63695 => x"ffffff",
   63696 => x"ffffff",
   63697 => x"ffffff",
   63698 => x"ffffff",
   63699 => x"ffffff",
   63700 => x"ffffff",
   63701 => x"ffffff",
   63702 => x"ffffff",
   63703 => x"ffffff",
   63704 => x"ffffff",
   63705 => x"ffffff",
   63706 => x"ffffff",
   63707 => x"ffffff",
   63708 => x"ffffff",
   63709 => x"ffffff",
   63710 => x"ffffff",
   63711 => x"ffffff",
   63712 => x"ffffff",
   63713 => x"ffffff",
   63714 => x"ffffff",
   63715 => x"ffffff",
   63716 => x"ffffff",
   63717 => x"ffffff",
   63718 => x"ffffff",
   63719 => x"ffffff",
   63720 => x"ffffff",
   63721 => x"ffffff",
   63722 => x"ffffff",
   63723 => x"ffffff",
   63724 => x"ffffff",
   63725 => x"ffffff",
   63726 => x"ffffff",
   63727 => x"ffffff",
   63728 => x"ffffff",
   63729 => x"ffffff",
   63730 => x"ffffff",
   63731 => x"ffffff",
   63732 => x"ffffff",
   63733 => x"ffffff",
   63734 => x"ffffff",
   63735 => x"ffffff",
   63736 => x"ffffff",
   63737 => x"ffffff",
   63738 => x"ffffff",
   63739 => x"ffffff",
   63740 => x"ffffff",
   63741 => x"ffffff",
   63742 => x"ffffff",
   63743 => x"ffffff",
   63744 => x"ffffff",
   63745 => x"ffffff",
   63746 => x"ffffff",
   63747 => x"ffffff",
   63748 => x"ffffff",
   63749 => x"ffffff",
   63750 => x"ffffff",
   63751 => x"ffffff",
   63752 => x"ffffff",
   63753 => x"ffffff",
   63754 => x"ffffff",
   63755 => x"ffffff",
   63756 => x"ffffff",
   63757 => x"ffffff",
   63758 => x"ffffff",
   63759 => x"ffffff",
   63760 => x"ffffff",
   63761 => x"ffffff",
   63762 => x"ffffff",
   63763 => x"ffffff",
   63764 => x"ffffff",
   63765 => x"ffffff",
   63766 => x"ffffff",
   63767 => x"ffffff",
   63768 => x"ffffff",
   63769 => x"ffffff",
   63770 => x"ffffff",
   63771 => x"ffffff",
   63772 => x"ffffff",
   63773 => x"ffffff",
   63774 => x"ffffff",
   63775 => x"ffffff",
   63776 => x"ffffff",
   63777 => x"ffffff",
   63778 => x"ffffff",
   63779 => x"ffffff",
   63780 => x"ffffff",
   63781 => x"ffffff",
   63782 => x"ffffff",
   63783 => x"ffffff",
   63784 => x"ffffff",
   63785 => x"ffffff",
   63786 => x"ffffff",
   63787 => x"ffffff",
   63788 => x"ffffff",
   63789 => x"ffffff",
   63790 => x"ffffff",
   63791 => x"ffffff",
   63792 => x"ffffff",
   63793 => x"ffffff",
   63794 => x"ffffff",
   63795 => x"ffffff",
   63796 => x"ffffff",
   63797 => x"ffffff",
   63798 => x"ffffff",
   63799 => x"ffffff",
   63800 => x"ffffff",
   63801 => x"ffffff",
   63802 => x"ffffff",
   63803 => x"ffffff",
   63804 => x"ffffff",
   63805 => x"ffffff",
   63806 => x"ffffff",
   63807 => x"ffffff",
   63808 => x"ffffff",
   63809 => x"ffffff",
   63810 => x"ffffff",
   63811 => x"ffffff",
   63812 => x"ffffff",
   63813 => x"ffffff",
   63814 => x"ffffff",
   63815 => x"ffffff",
   63816 => x"ffffff",
   63817 => x"ffffff",
   63818 => x"ffffff",
   63819 => x"ffffff",
   63820 => x"ffffff",
   63821 => x"ffffff",
   63822 => x"ffffff",
   63823 => x"ffffff",
   63824 => x"ffffff",
   63825 => x"ffffff",
   63826 => x"ffffff",
   63827 => x"ffffff",
   63828 => x"ffffff",
   63829 => x"ffffff",
   63830 => x"ffffff",
   63831 => x"ffffff",
   63832 => x"ffffff",
   63833 => x"ffffff",
   63834 => x"ffffff",
   63835 => x"ffffff",
   63836 => x"ffffff",
   63837 => x"ffffff",
   63838 => x"ffffff",
   63839 => x"ffffff",
   63840 => x"ffffff",
   63841 => x"ffffff",
   63842 => x"ffffff",
   63843 => x"ffffff",
   63844 => x"ffffff",
   63845 => x"ffffff",
   63846 => x"ffffff",
   63847 => x"ffffff",
   63848 => x"ffffff",
   63849 => x"ffffff",
   63850 => x"ffffff",
   63851 => x"ffffff",
   63852 => x"ffffff",
   63853 => x"ffffff",
   63854 => x"ffffff",
   63855 => x"ffffff",
   63856 => x"ffffff",
   63857 => x"ffffff",
   63858 => x"ffffff",
   63859 => x"ffffff",
   63860 => x"ffffff",
   63861 => x"ffffff",
   63862 => x"ffffff",
   63863 => x"ffffff",
   63864 => x"ffffff",
   63865 => x"ffffff",
   63866 => x"ffffff",
   63867 => x"ffffff",
   63868 => x"ffffff",
   63869 => x"ffffff",
   63870 => x"ffffff",
   63871 => x"ffffff",
   63872 => x"ffffff",
   63873 => x"ffffff",
   63874 => x"ffffff",
   63875 => x"ffffff",
   63876 => x"ffffff",
   63877 => x"ffffff",
   63878 => x"ffffff",
   63879 => x"ffffff",
   63880 => x"ffffff",
   63881 => x"ffffff",
   63882 => x"ffffff",
   63883 => x"ffffff",
   63884 => x"ffffff",
   63885 => x"ffffff",
   63886 => x"ffffff",
   63887 => x"ffffff",
   63888 => x"ffffff",
   63889 => x"ffffff",
   63890 => x"ffffff",
   63891 => x"ffffff",
   63892 => x"ffffff",
   63893 => x"ffffff",
   63894 => x"ffffff",
   63895 => x"ffffff",
   63896 => x"ffffff",
   63897 => x"ffffff",
   63898 => x"ffffff",
   63899 => x"ffffff",
   63900 => x"ffffff",
   63901 => x"ffffff",
   63902 => x"ffffff",
   63903 => x"ffffff",
   63904 => x"ffffff",
   63905 => x"ffffff",
   63906 => x"ffffff",
   63907 => x"ffffff",
   63908 => x"ffffff",
   63909 => x"ffffff",
   63910 => x"ffffff",
   63911 => x"ffffff",
   63912 => x"ffffff",
   63913 => x"ffffff",
   63914 => x"ffffff",
   63915 => x"ffffff",
   63916 => x"ffffff",
   63917 => x"ffffff",
   63918 => x"ffffff",
   63919 => x"ffffff",
   63920 => x"ffffff",
   63921 => x"ffffff",
   63922 => x"ffffff",
   63923 => x"ffffff",
   63924 => x"ffffff",
   63925 => x"ffffff",
   63926 => x"ffffff",
   63927 => x"ffffff",
   63928 => x"ffffff",
   63929 => x"ffffff",
   63930 => x"ffffff",
   63931 => x"ffffff",
   63932 => x"ffffff",
   63933 => x"ffffff",
   63934 => x"ffffff",
   63935 => x"ffffff",
   63936 => x"ffffff",
   63937 => x"ffffff",
   63938 => x"ffffff",
   63939 => x"ffffff",
   63940 => x"ffffff",
   63941 => x"ffffff",
   63942 => x"ffffff",
   63943 => x"ffffff",
   63944 => x"ffffff",
   63945 => x"ffffff",
   63946 => x"ffffff",
   63947 => x"ffffff",
   63948 => x"ffffff",
   63949 => x"ffffff",
   63950 => x"ffffff",
   63951 => x"ffffff",
   63952 => x"ffffff",
   63953 => x"ffffff",
   63954 => x"ffffff",
   63955 => x"ffffff",
   63956 => x"ffffff",
   63957 => x"ffffff",
   63958 => x"ffffff",
   63959 => x"ffffff",
   63960 => x"ffffff",
   63961 => x"ffffff",
   63962 => x"ffffff",
   63963 => x"ffffff",
   63964 => x"ffffff",
   63965 => x"ffffff",
   63966 => x"ffffff",
   63967 => x"ffffff",
   63968 => x"ffffff",
   63969 => x"ffffff",
   63970 => x"ffffff",
   63971 => x"ffffff",
   63972 => x"ffffff",
   63973 => x"ffffff",
   63974 => x"ffffff",
   63975 => x"ffffff",
   63976 => x"ffffff",
   63977 => x"ffffff",
   63978 => x"ffffff",
   63979 => x"ffffff",
   63980 => x"ffffff",
   63981 => x"ffffff",
   63982 => x"ffffff",
   63983 => x"ffffff",
   63984 => x"ffffff",
   63985 => x"ffffff",
   63986 => x"ffffff",
   63987 => x"ffffff",
   63988 => x"ffffff",
   63989 => x"ffffff",
   63990 => x"ffffff",
   63991 => x"ffffff",
   63992 => x"ffffff",
   63993 => x"ffffff",
   63994 => x"ffffff",
   63995 => x"ffffff",
   63996 => x"ffffff",
   63997 => x"ffffff",
   63998 => x"ffffff",
   63999 => x"ffffff",
   64000 => x"ffffff",
   64001 => x"ffffff",
   64002 => x"ffffff",
   64003 => x"ffffff",
   64004 => x"ffffff",
   64005 => x"ffffff",
   64006 => x"ffffff",
   64007 => x"ffffff",
   64008 => x"ffffff",
   64009 => x"ffffff",
   64010 => x"ffffff",
   64011 => x"ffffff",
   64012 => x"ffffff",
   64013 => x"ffffff",
   64014 => x"ffffff",
   64015 => x"ffffff",
   64016 => x"ffffff",
   64017 => x"ffffff",
   64018 => x"ffffff",
   64019 => x"ffffff",
   64020 => x"ffffff",
   64021 => x"ffffff",
   64022 => x"ffffff",
   64023 => x"ffffff",
   64024 => x"ffffff",
   64025 => x"ffffff",
   64026 => x"ffffff",
   64027 => x"ffffff",
   64028 => x"ffffff",
   64029 => x"ffffff",
   64030 => x"ffffff",
   64031 => x"ffffff",
   64032 => x"ffffff",
   64033 => x"ffffff",
   64034 => x"ffffff",
   64035 => x"ffffff",
   64036 => x"ffffff",
   64037 => x"ffffff",
   64038 => x"ffffff",
   64039 => x"ffffff",
   64040 => x"ffffff",
   64041 => x"ffffff",
   64042 => x"ffffff",
   64043 => x"ffffff",
   64044 => x"ffffff",
   64045 => x"ffffff",
   64046 => x"ffffff",
   64047 => x"ffffff",
   64048 => x"ffffff",
   64049 => x"ffffff",
   64050 => x"ffffff",
   64051 => x"ffffff",
   64052 => x"ffffff",
   64053 => x"ffffff",
   64054 => x"ffffff",
   64055 => x"ffffff",
   64056 => x"ffffff",
   64057 => x"ffffff",
   64058 => x"ffffff",
   64059 => x"ffffff",
   64060 => x"ffffff",
   64061 => x"ffffff",
   64062 => x"ffffff",
   64063 => x"ffffff",
   64064 => x"ffffff",
   64065 => x"ffffff",
   64066 => x"ffffff",
   64067 => x"ffffff",
   64068 => x"ffffff",
   64069 => x"ffffff",
   64070 => x"ffffff",
   64071 => x"ffffff",
   64072 => x"ffffff",
   64073 => x"ffffff",
   64074 => x"ffffff",
   64075 => x"ffffff",
   64076 => x"ffffff",
   64077 => x"ffffff",
   64078 => x"ffffff",
   64079 => x"ffffff",
   64080 => x"ffffff",
   64081 => x"ffffff",
   64082 => x"ffffff",
   64083 => x"ffffff",
   64084 => x"ffffff",
   64085 => x"ffffff",
   64086 => x"ffffff",
   64087 => x"ffffff",
   64088 => x"ffffff",
   64089 => x"ffffff",
   64090 => x"ffffff",
   64091 => x"ffffff",
   64092 => x"ffffff",
   64093 => x"ffffff",
   64094 => x"ffffff",
   64095 => x"ffffff",
   64096 => x"ffffff",
   64097 => x"ffffff",
   64098 => x"ffffff",
   64099 => x"ffffff",
   64100 => x"ffffff",
   64101 => x"ffffff",
   64102 => x"ffffff",
   64103 => x"ffffff",
   64104 => x"ffffff",
   64105 => x"ffffff",
   64106 => x"ffffff",
   64107 => x"ffffff",
   64108 => x"ffffff",
   64109 => x"ffffff",
   64110 => x"ffffff",
   64111 => x"ffffff",
   64112 => x"ffffff",
   64113 => x"ffffff",
   64114 => x"ffffff",
   64115 => x"ffffff",
   64116 => x"ffffff",
   64117 => x"ffffff",
   64118 => x"ffffff",
   64119 => x"ffffff",
   64120 => x"ffffff",
   64121 => x"ffffff",
   64122 => x"ffffff",
   64123 => x"ffffff",
   64124 => x"ffffff",
   64125 => x"ffffff",
   64126 => x"ffffff",
   64127 => x"ffffff",
   64128 => x"ffffff",
   64129 => x"ffffff",
   64130 => x"ffffff",
   64131 => x"ffffff",
   64132 => x"ffffff",
   64133 => x"ffffff",
   64134 => x"ffffff",
   64135 => x"ffffff",
   64136 => x"ffffff",
   64137 => x"ffffff",
   64138 => x"ffffff",
   64139 => x"ffffff",
   64140 => x"ffffff",
   64141 => x"ffffff",
   64142 => x"ffffff",
   64143 => x"ffffff",
   64144 => x"ffffff",
   64145 => x"ffffff",
   64146 => x"ffffff",
   64147 => x"ffffff",
   64148 => x"ffffff",
   64149 => x"ffffff",
   64150 => x"ffffff",
   64151 => x"ffffff",
   64152 => x"ffffff",
   64153 => x"ffffff",
   64154 => x"ffffff",
   64155 => x"ffffff",
   64156 => x"ffffff",
   64157 => x"ffffff",
   64158 => x"ffffff",
   64159 => x"ffffff",
   64160 => x"ffffff",
   64161 => x"ffffff",
   64162 => x"ffffff",
   64163 => x"ffffff",
   64164 => x"ffffff",
   64165 => x"ffffff",
   64166 => x"ffffff",
   64167 => x"ffffff",
   64168 => x"ffffff",
   64169 => x"ffffff",
   64170 => x"ffffff",
   64171 => x"ffffff",
   64172 => x"ffffff",
   64173 => x"ffffff",
   64174 => x"ffffff",
   64175 => x"ffffff",
   64176 => x"ffffff",
   64177 => x"ffffff",
   64178 => x"ffffff",
   64179 => x"ffffff",
   64180 => x"ffffff",
   64181 => x"ffffff",
   64182 => x"ffffff",
   64183 => x"ffffff",
   64184 => x"ffffff",
   64185 => x"ffffff",
   64186 => x"ffffff",
   64187 => x"ffffff",
   64188 => x"ffffff",
   64189 => x"ffffff",
   64190 => x"ffffff",
   64191 => x"ffffff",
   64192 => x"ffffff",
   64193 => x"ffffff",
   64194 => x"ffffff",
   64195 => x"ffffff",
   64196 => x"ffffff",
   64197 => x"ffffff",
   64198 => x"ffffff",
   64199 => x"ffffff",
   64200 => x"ffffff",
   64201 => x"ffffff",
   64202 => x"ffffff",
   64203 => x"ffffff",
   64204 => x"ffffff",
   64205 => x"ffffff",
   64206 => x"ffffff",
   64207 => x"ffffff",
   64208 => x"ffffff",
   64209 => x"ffffff",
   64210 => x"ffffff",
   64211 => x"ffffff",
   64212 => x"ffffff",
   64213 => x"ffffff",
   64214 => x"ffffff",
   64215 => x"ffffff",
   64216 => x"ffffff",
   64217 => x"ffffff",
   64218 => x"ffffff",
   64219 => x"ffffff",
   64220 => x"ffffff",
   64221 => x"ffffff",
   64222 => x"ffffff",
   64223 => x"ffffff",
   64224 => x"ffffff",
   64225 => x"ffffff",
   64226 => x"ffffff",
   64227 => x"ffffff",
   64228 => x"ffffff",
   64229 => x"ffffff",
   64230 => x"ffffff",
   64231 => x"ffffff",
   64232 => x"ffffff",
   64233 => x"ffffff",
   64234 => x"ffffff",
   64235 => x"ffffff",
   64236 => x"ffffff",
   64237 => x"ffffff",
   64238 => x"ffffff",
   64239 => x"ffffff",
   64240 => x"ffffff",
   64241 => x"ffffff",
   64242 => x"ffffff",
   64243 => x"ffffff",
   64244 => x"ffffff",
   64245 => x"ffffff",
   64246 => x"ffffff",
   64247 => x"ffffff",
   64248 => x"ffffff",
   64249 => x"ffffff",
   64250 => x"ffffff",
   64251 => x"ffffff",
   64252 => x"ffffff",
   64253 => x"ffffff",
   64254 => x"ffffff",
   64255 => x"ffffff",
   64256 => x"ffffff",
   64257 => x"ffffff",
   64258 => x"ffffff",
   64259 => x"ffffff",
   64260 => x"ffffff",
   64261 => x"ffffff",
   64262 => x"ffffff",
   64263 => x"ffffff",
   64264 => x"ffffff",
   64265 => x"ffffff",
   64266 => x"ffffff",
   64267 => x"ffffff",
   64268 => x"ffffff",
   64269 => x"ffffff",
   64270 => x"ffffff",
   64271 => x"ffffff",
   64272 => x"ffffff",
   64273 => x"ffffff",
   64274 => x"ffffff",
   64275 => x"ffffff",
   64276 => x"ffffff",
   64277 => x"ffffff",
   64278 => x"ffffff",
   64279 => x"ffffff",
   64280 => x"ffffff",
   64281 => x"ffffff",
   64282 => x"ffffff",
   64283 => x"ffffff",
   64284 => x"ffffff",
   64285 => x"ffffff",
   64286 => x"ffffff",
   64287 => x"ffffff",
   64288 => x"ffffff",
   64289 => x"ffffff",
   64290 => x"ffffff",
   64291 => x"ffffff",
   64292 => x"ffffff",
   64293 => x"ffffff",
   64294 => x"ffffff",
   64295 => x"ffffff",
   64296 => x"ffffff",
   64297 => x"ffffff",
   64298 => x"ffffff",
   64299 => x"ffffff",
   64300 => x"ffffff",
   64301 => x"ffffff",
   64302 => x"ffffff",
   64303 => x"ffffff",
   64304 => x"ffffff",
   64305 => x"ffffff",
   64306 => x"ffffff",
   64307 => x"ffffff",
   64308 => x"ffffff",
   64309 => x"ffffff",
   64310 => x"ffffff",
   64311 => x"ffffff",
   64312 => x"ffffff",
   64313 => x"ffffff",
   64314 => x"ffffff",
   64315 => x"ffffff",
   64316 => x"ffffff",
   64317 => x"ffffff",
   64318 => x"ffffff",
   64319 => x"ffffff",
   64320 => x"ffffff",
   64321 => x"ffffff",
   64322 => x"ffffff",
   64323 => x"ffffff",
   64324 => x"ffffff",
   64325 => x"ffffff",
   64326 => x"ffffff",
   64327 => x"ffffff",
   64328 => x"ffffff",
   64329 => x"ffffff",
   64330 => x"ffffff",
   64331 => x"ffffff",
   64332 => x"ffffff",
   64333 => x"ffffff",
   64334 => x"ffffff",
   64335 => x"ffffff",
   64336 => x"ffffff",
   64337 => x"ffffff",
   64338 => x"ffffff",
   64339 => x"ffffff",
   64340 => x"ffffff",
   64341 => x"ffffff",
   64342 => x"ffffff",
   64343 => x"ffffff",
   64344 => x"ffffff",
   64345 => x"ffffff",
   64346 => x"ffffff",
   64347 => x"ffffff",
   64348 => x"ffffff",
   64349 => x"ffffff",
   64350 => x"ffffff",
   64351 => x"ffffff",
   64352 => x"ffffff",
   64353 => x"ffffff",
   64354 => x"ffffff",
   64355 => x"ffffff",
   64356 => x"ffffff",
   64357 => x"ffffff",
   64358 => x"ffffff",
   64359 => x"ffffff",
   64360 => x"ffffff",
   64361 => x"ffffff",
   64362 => x"ffffff",
   64363 => x"ffffff",
   64364 => x"ffffff",
   64365 => x"ffffff",
   64366 => x"ffffff",
   64367 => x"ffffff",
   64368 => x"ffffff",
   64369 => x"ffffff",
   64370 => x"ffffff",
   64371 => x"ffffff",
   64372 => x"ffffff",
   64373 => x"ffffff",
   64374 => x"ffffff",
   64375 => x"ffffff",
   64376 => x"ffffff",
   64377 => x"ffffff",
   64378 => x"ffffff",
   64379 => x"ffffff",
   64380 => x"ffffff",
   64381 => x"ffffff",
   64382 => x"ffffff",
   64383 => x"ffffff",
   64384 => x"ffffff",
   64385 => x"ffffff",
   64386 => x"ffffff",
   64387 => x"ffffff",
   64388 => x"ffffff",
   64389 => x"ffffff",
   64390 => x"ffffff",
   64391 => x"ffffff",
   64392 => x"ffffff",
   64393 => x"ffffff",
   64394 => x"ffffff",
   64395 => x"ffffff",
   64396 => x"ffffff",
   64397 => x"ffffff",
   64398 => x"ffffff",
   64399 => x"ffffff",
   64400 => x"ffffff",
   64401 => x"ffffff",
   64402 => x"ffffff",
   64403 => x"ffffff",
   64404 => x"ffffff",
   64405 => x"ffffff",
   64406 => x"ffffff",
   64407 => x"ffffff",
   64408 => x"ffffff",
   64409 => x"ffffff",
   64410 => x"ffffff",
   64411 => x"ffffff",
   64412 => x"ffffff",
   64413 => x"ffffff",
   64414 => x"ffffff",
   64415 => x"ffffff",
   64416 => x"ffffff",
   64417 => x"ffffff",
   64418 => x"ffffff",
   64419 => x"ffffff",
   64420 => x"ffffff",
   64421 => x"ffffff",
   64422 => x"ffffff",
   64423 => x"ffffff",
   64424 => x"ffffff",
   64425 => x"ffffff",
   64426 => x"ffffff",
   64427 => x"ffffff",
   64428 => x"ffffff",
   64429 => x"ffffff",
   64430 => x"ffffff",
   64431 => x"ffffff",
   64432 => x"ffffff",
   64433 => x"ffffff",
   64434 => x"ffffff",
   64435 => x"ffffff",
   64436 => x"ffffff",
   64437 => x"ffffff",
   64438 => x"ffffff",
   64439 => x"ffffff",
   64440 => x"ffffff",
   64441 => x"ffffff",
   64442 => x"ffffff",
   64443 => x"ffffff",
   64444 => x"ffffff",
   64445 => x"ffffff",
   64446 => x"ffffff",
   64447 => x"ffffff",
   64448 => x"ffffff",
   64449 => x"ffffff",
   64450 => x"ffffff",
   64451 => x"ffffff",
   64452 => x"ffffff",
   64453 => x"ffffff",
   64454 => x"ffffff",
   64455 => x"ffffff",
   64456 => x"ffffff",
   64457 => x"ffffff",
   64458 => x"ffffff",
   64459 => x"ffffff",
   64460 => x"ffffff",
   64461 => x"ffffff",
   64462 => x"ffffff",
   64463 => x"ffffff",
   64464 => x"ffffff",
   64465 => x"ffffff",
   64466 => x"ffffff",
   64467 => x"ffffff",
   64468 => x"ffffff",
   64469 => x"ffffff",
   64470 => x"ffffff",
   64471 => x"ffffff",
   64472 => x"ffffff",
   64473 => x"ffffff",
   64474 => x"ffffff",
   64475 => x"ffffff",
   64476 => x"ffffff",
   64477 => x"ffffff",
   64478 => x"ffffff",
   64479 => x"ffffff",
   64480 => x"ffffff",
   64481 => x"ffffff",
   64482 => x"ffffff",
   64483 => x"ffffff",
   64484 => x"ffffff",
   64485 => x"ffffff",
   64486 => x"ffffff",
   64487 => x"ffffff",
   64488 => x"ffffff",
   64489 => x"ffffff",
   64490 => x"ffffff",
   64491 => x"ffffff",
   64492 => x"ffffff",
   64493 => x"ffffff",
   64494 => x"ffffff",
   64495 => x"ffffff",
   64496 => x"ffffff",
   64497 => x"ffffff",
   64498 => x"ffffff",
   64499 => x"ffffff",
   64500 => x"ffffff",
   64501 => x"ffffff",
   64502 => x"ffffff",
   64503 => x"ffffff",
   64504 => x"ffffff",
   64505 => x"ffffff",
   64506 => x"ffffff",
   64507 => x"ffffff",
   64508 => x"ffffff",
   64509 => x"ffffff",
   64510 => x"ffffff",
   64511 => x"ffffff",
   64512 => x"ffffff",
   64513 => x"ffffff",
   64514 => x"ffffff",
   64515 => x"ffffff",
   64516 => x"ffffff",
   64517 => x"ffffff",
   64518 => x"ffffff",
   64519 => x"ffffff",
   64520 => x"ffffff",
   64521 => x"ffffff",
   64522 => x"ffffff",
   64523 => x"ffffff",
   64524 => x"ffffff",
   64525 => x"ffffff",
   64526 => x"ffffff",
   64527 => x"ffffff",
   64528 => x"ffffff",
   64529 => x"ffffff",
   64530 => x"ffffff",
   64531 => x"ffffff",
   64532 => x"ffffff",
   64533 => x"ffffff",
   64534 => x"ffffff",
   64535 => x"ffffff",
   64536 => x"ffffff",
   64537 => x"ffffff",
   64538 => x"ffffff",
   64539 => x"ffffff",
   64540 => x"ffffff",
   64541 => x"ffffff",
   64542 => x"ffffff",
   64543 => x"ffffff",
   64544 => x"ffffff",
   64545 => x"ffffff",
   64546 => x"ffffff",
   64547 => x"ffffff",
   64548 => x"ffffff",
   64549 => x"ffffff",
   64550 => x"ffffff",
   64551 => x"ffffff",
   64552 => x"ffffff",
   64553 => x"ffffff",
   64554 => x"ffffff",
   64555 => x"ffffff",
   64556 => x"ffffff",
   64557 => x"ffffff",
   64558 => x"ffffff",
   64559 => x"ffffff",
   64560 => x"ffffff",
   64561 => x"ffffff",
   64562 => x"ffffff",
   64563 => x"ffffff",
   64564 => x"ffffff",
   64565 => x"ffffff",
   64566 => x"ffffff",
   64567 => x"ffffff",
   64568 => x"ffffff",
   64569 => x"ffffff",
   64570 => x"ffffff",
   64571 => x"ffffff",
   64572 => x"ffffff",
   64573 => x"ffffff",
   64574 => x"ffffff",
   64575 => x"ffffff",
   64576 => x"ffffff",
   64577 => x"ffffff",
   64578 => x"ffffff",
   64579 => x"ffffff",
   64580 => x"ffffff",
   64581 => x"ffffff",
   64582 => x"ffffff",
   64583 => x"ffffff",
   64584 => x"ffffff",
   64585 => x"ffffff",
   64586 => x"ffffff",
   64587 => x"ffffff",
   64588 => x"ffffff",
   64589 => x"ffffff",
   64590 => x"ffffff",
   64591 => x"ffffff",
   64592 => x"ffffff",
   64593 => x"ffffff",
   64594 => x"ffffff",
   64595 => x"ffffff",
   64596 => x"ffffff",
   64597 => x"ffffff",
   64598 => x"ffffff",
   64599 => x"ffffff",
   64600 => x"ffffff",
   64601 => x"ffffff",
   64602 => x"ffffff",
   64603 => x"ffffff",
   64604 => x"ffffff",
   64605 => x"ffffff",
   64606 => x"ffffff",
   64607 => x"ffffff",
   64608 => x"ffffff",
   64609 => x"ffffff",
   64610 => x"ffffff",
   64611 => x"ffffff",
   64612 => x"ffffff",
   64613 => x"ffffff",
   64614 => x"ffffff",
   64615 => x"ffffff",
   64616 => x"ffffff",
   64617 => x"ffffff",
   64618 => x"ffffff",
   64619 => x"ffffff",
   64620 => x"ffffff",
   64621 => x"ffffff",
   64622 => x"ffffff",
   64623 => x"ffffff",
   64624 => x"ffffff",
   64625 => x"ffffff",
   64626 => x"ffffff",
   64627 => x"ffffff",
   64628 => x"ffffff",
   64629 => x"ffffff",
   64630 => x"ffffff",
   64631 => x"ffffff",
   64632 => x"ffffff",
   64633 => x"ffffff",
   64634 => x"ffffff",
   64635 => x"ffffff",
   64636 => x"ffffff",
   64637 => x"ffffff",
   64638 => x"ffffff",
   64639 => x"ffffff",
   64640 => x"ffffff",
   64641 => x"ffffff",
   64642 => x"ffffff",
   64643 => x"ffffff",
   64644 => x"ffffff",
   64645 => x"ffffff",
   64646 => x"ffffff",
   64647 => x"ffffff",
   64648 => x"ffffff",
   64649 => x"ffffff",
   64650 => x"ffffff",
   64651 => x"ffffff",
   64652 => x"ffffff",
   64653 => x"ffffff",
   64654 => x"ffffff",
   64655 => x"ffffff",
   64656 => x"ffffff",
   64657 => x"ffffff",
   64658 => x"ffffff",
   64659 => x"ffffff",
   64660 => x"ffffff",
   64661 => x"ffffff",
   64662 => x"ffffff",
   64663 => x"ffffff",
   64664 => x"ffffff",
   64665 => x"ffffff",
   64666 => x"ffffff",
   64667 => x"ffffff",
   64668 => x"ffffff",
   64669 => x"ffffff",
   64670 => x"ffffff",
   64671 => x"ffffff",
   64672 => x"ffffff",
   64673 => x"ffffff",
   64674 => x"ffffff",
   64675 => x"ffffff",
   64676 => x"ffffff",
   64677 => x"ffffff",
   64678 => x"ffffff",
   64679 => x"ffffff",
   64680 => x"ffffff",
   64681 => x"ffffff",
   64682 => x"ffffff",
   64683 => x"ffffff",
   64684 => x"ffffff",
   64685 => x"ffffff",
   64686 => x"ffffff",
   64687 => x"ffffff",
   64688 => x"ffffff",
   64689 => x"ffffff",
   64690 => x"ffffff",
   64691 => x"ffffff",
   64692 => x"ffffff",
   64693 => x"ffffff",
   64694 => x"ffffff",
   64695 => x"ffffff",
   64696 => x"ffffff",
   64697 => x"ffffff",
   64698 => x"ffffff",
   64699 => x"ffffff",
   64700 => x"ffffff",
   64701 => x"ffffff",
   64702 => x"ffffff",
   64703 => x"ffffff",
   64704 => x"ffffff",
   64705 => x"ffffff",
   64706 => x"ffffff",
   64707 => x"ffffff",
   64708 => x"ffffff",
   64709 => x"ffffff",
   64710 => x"ffffff",
   64711 => x"ffffff",
   64712 => x"ffffff",
   64713 => x"ffffff",
   64714 => x"ffffff",
   64715 => x"ffffff",
   64716 => x"ffffff",
   64717 => x"ffffff",
   64718 => x"ffffff",
   64719 => x"ffffff",
   64720 => x"ffffff",
   64721 => x"ffffff",
   64722 => x"ffffff",
   64723 => x"ffffff",
   64724 => x"ffffff",
   64725 => x"ffffff",
   64726 => x"ffffff",
   64727 => x"ffffff",
   64728 => x"ffffff",
   64729 => x"ffffff",
   64730 => x"ffffff",
   64731 => x"ffffff",
   64732 => x"ffffff",
   64733 => x"ffffff",
   64734 => x"ffffff",
   64735 => x"ffffff",
   64736 => x"ffffff",
   64737 => x"ffffff",
   64738 => x"ffffff",
   64739 => x"ffffff",
   64740 => x"ffffff",
   64741 => x"ffffff",
   64742 => x"ffffff",
   64743 => x"ffffff",
   64744 => x"ffffff",
   64745 => x"ffffff",
   64746 => x"ffffff",
   64747 => x"ffffff",
   64748 => x"ffffff",
   64749 => x"ffffff",
   64750 => x"ffffff",
   64751 => x"ffffff",
   64752 => x"ffffff",
   64753 => x"ffffff",
   64754 => x"ffffff",
   64755 => x"ffffff",
   64756 => x"ffffff",
   64757 => x"ffffff",
   64758 => x"ffffff",
   64759 => x"ffffff",
   64760 => x"ffffff",
   64761 => x"ffffff",
   64762 => x"ffffff",
   64763 => x"ffffff",
   64764 => x"ffffff",
   64765 => x"ffffff",
   64766 => x"ffffff",
   64767 => x"ffffff",
   64768 => x"ffffff",
   64769 => x"ffffff",
   64770 => x"ffffff",
   64771 => x"ffffff",
   64772 => x"ffffff",
   64773 => x"ffffff",
   64774 => x"ffffff",
   64775 => x"ffffff",
   64776 => x"ffffff",
   64777 => x"ffffff",
   64778 => x"ffffff",
   64779 => x"ffffff",
   64780 => x"ffffff",
   64781 => x"ffffff",
   64782 => x"ffffff",
   64783 => x"ffffff",
   64784 => x"ffffff",
   64785 => x"ffffff",
   64786 => x"ffffff",
   64787 => x"ffffff",
   64788 => x"ffffff",
   64789 => x"ffffff",
   64790 => x"ffffff",
   64791 => x"ffffff",
   64792 => x"ffffff",
   64793 => x"ffffff",
   64794 => x"ffffff",
   64795 => x"ffffff",
   64796 => x"ffffff",
   64797 => x"ffffff",
   64798 => x"ffffff",
   64799 => x"ffffff",
   64800 => x"ffffff",
   64801 => x"ffffff",
   64802 => x"ffffff",
   64803 => x"ffffff",
   64804 => x"ffffff",
   64805 => x"ffffff",
   64806 => x"ffffff",
   64807 => x"ffffff",
   64808 => x"ffffff",
   64809 => x"ffffff",
   64810 => x"ffffff",
   64811 => x"ffffff",
   64812 => x"ffffff",
   64813 => x"ffffff",
   64814 => x"ffffff",
   64815 => x"ffffff",
   64816 => x"ffffff",
   64817 => x"ffffff",
   64818 => x"ffffff",
   64819 => x"ffffff",
   64820 => x"ffffff",
   64821 => x"ffffff",
   64822 => x"ffffff",
   64823 => x"ffffff",
   64824 => x"ffffff",
   64825 => x"ffffff",
   64826 => x"ffffff",
   64827 => x"ffffff",
   64828 => x"ffffff",
   64829 => x"ffffff",
   64830 => x"ffffff",
   64831 => x"ffffff",
   64832 => x"ffffff",
   64833 => x"ffffff",
   64834 => x"ffffff",
   64835 => x"ffffff",
   64836 => x"ffffff",
   64837 => x"ffffff",
   64838 => x"ffffff",
   64839 => x"ffffff",
   64840 => x"ffffff",
   64841 => x"ffffff",
   64842 => x"ffffff",
   64843 => x"ffffff",
   64844 => x"ffffff",
   64845 => x"ffffff",
   64846 => x"ffffff",
   64847 => x"ffffff",
   64848 => x"ffffff",
   64849 => x"ffffff",
   64850 => x"ffffff",
   64851 => x"ffffff",
   64852 => x"ffffff",
   64853 => x"ffffff",
   64854 => x"ffffff",
   64855 => x"ffffff",
   64856 => x"ffffff",
   64857 => x"ffffff",
   64858 => x"ffffff",
   64859 => x"ffffff",
   64860 => x"ffffff",
   64861 => x"ffffff",
   64862 => x"ffffff",
   64863 => x"ffffff",
   64864 => x"ffffff",
   64865 => x"ffffff",
   64866 => x"ffffff",
   64867 => x"ffffff",
   64868 => x"ffffff",
   64869 => x"ffffff",
   64870 => x"ffffff",
   64871 => x"ffffff",
   64872 => x"ffffff",
   64873 => x"ffffff",
   64874 => x"ffffff",
   64875 => x"ffffff",
   64876 => x"ffffff",
   64877 => x"ffffff",
   64878 => x"ffffff",
   64879 => x"ffffff",
   64880 => x"ffffff",
   64881 => x"ffffff",
   64882 => x"ffffff",
   64883 => x"ffffff",
   64884 => x"ffffff",
   64885 => x"ffffff",
   64886 => x"ffffff",
   64887 => x"ffffff",
   64888 => x"ffffff",
   64889 => x"ffffff",
   64890 => x"ffffff",
   64891 => x"ffffff",
   64892 => x"ffffff",
   64893 => x"ffffff",
   64894 => x"ffffff",
   64895 => x"ffffff",
   64896 => x"ffffff",
   64897 => x"ffffff",
   64898 => x"ffffff",
   64899 => x"ffffff",
   64900 => x"ffffff",
   64901 => x"ffffff",
   64902 => x"ffffff",
   64903 => x"ffffff",
   64904 => x"ffffff",
   64905 => x"ffffff",
   64906 => x"ffffff",
   64907 => x"ffffff",
   64908 => x"ffffff",
   64909 => x"ffffff",
   64910 => x"ffffff",
   64911 => x"ffffff",
   64912 => x"ffffff",
   64913 => x"ffffff",
   64914 => x"ffffff",
   64915 => x"ffffff",
   64916 => x"ffffff",
   64917 => x"ffffff",
   64918 => x"ffffff",
   64919 => x"ffffff",
   64920 => x"ffffff",
   64921 => x"ffffff",
   64922 => x"ffffff",
   64923 => x"ffffff",
   64924 => x"ffffff",
   64925 => x"ffffff",
   64926 => x"ffffff",
   64927 => x"ffffff",
   64928 => x"ffffff",
   64929 => x"ffffff",
   64930 => x"ffffff",
   64931 => x"ffffff",
   64932 => x"ffffff",
   64933 => x"ffffff",
   64934 => x"ffffff",
   64935 => x"ffffff",
   64936 => x"ffffff",
   64937 => x"ffffff",
   64938 => x"ffffff",
   64939 => x"ffffff",
   64940 => x"ffffff",
   64941 => x"ffffff",
   64942 => x"ffffff",
   64943 => x"ffffff",
   64944 => x"ffffff",
   64945 => x"ffffff",
   64946 => x"ffffff",
   64947 => x"ffffff",
   64948 => x"ffffff",
   64949 => x"ffffff",
   64950 => x"ffffff",
   64951 => x"ffffff",
   64952 => x"ffffff",
   64953 => x"ffffff",
   64954 => x"ffffff",
   64955 => x"ffffff",
   64956 => x"ffffff",
   64957 => x"ffffff",
   64958 => x"ffffff",
   64959 => x"ffffff",
   64960 => x"ffffff",
   64961 => x"ffffff",
   64962 => x"ffffff",
   64963 => x"ffffff",
   64964 => x"ffffff",
   64965 => x"ffffff",
   64966 => x"ffffff",
   64967 => x"ffffff",
   64968 => x"ffffff",
   64969 => x"ffffff",
   64970 => x"ffffff",
   64971 => x"ffffff",
   64972 => x"ffffff",
   64973 => x"ffffff",
   64974 => x"ffffff",
   64975 => x"ffffff",
   64976 => x"ffffff",
   64977 => x"ffffff",
   64978 => x"ffffff",
   64979 => x"ffffff",
   64980 => x"ffffff",
   64981 => x"ffffff",
   64982 => x"ffffff",
   64983 => x"ffffff",
   64984 => x"ffffff",
   64985 => x"ffffff",
   64986 => x"ffffff",
   64987 => x"ffffff",
   64988 => x"ffffff",
   64989 => x"ffffff",
   64990 => x"ffffff",
   64991 => x"ffffff",
   64992 => x"ffffff",
   64993 => x"ffffff",
   64994 => x"ffffff",
   64995 => x"ffffff",
   64996 => x"ffffff",
   64997 => x"ffffff",
   64998 => x"ffffff",
   64999 => x"ffffff",
   65000 => x"ffffff",
   65001 => x"ffffff",
   65002 => x"ffffff",
   65003 => x"ffffff",
   65004 => x"ffffff",
   65005 => x"ffffff",
   65006 => x"ffffff",
   65007 => x"ffffff",
   65008 => x"ffffff",
   65009 => x"ffffff",
   65010 => x"ffffff",
   65011 => x"ffffff",
   65012 => x"ffffff",
   65013 => x"ffffff",
   65014 => x"ffffff",
   65015 => x"ffffff",
   65016 => x"ffffff",
   65017 => x"ffffff",
   65018 => x"ffffff",
   65019 => x"ffffff",
   65020 => x"ffffff",
   65021 => x"ffffff",
   65022 => x"ffffff",
   65023 => x"ffffff",
   65024 => x"ffffff",
   65025 => x"ffffff",
   65026 => x"ffffff",
   65027 => x"ffffff",
   65028 => x"ffffff",
   65029 => x"ffffff",
   65030 => x"ffffff",
   65031 => x"ffffff",
   65032 => x"ffffff",
   65033 => x"ffffff",
   65034 => x"ffffff",
   65035 => x"ffffff",
   65036 => x"ffffff",
   65037 => x"ffffff",
   65038 => x"ffffff",
   65039 => x"ffffff",
   65040 => x"ffffff",
   65041 => x"ffffff",
   65042 => x"ffffff",
   65043 => x"ffffff",
   65044 => x"ffffff",
   65045 => x"ffffff",
   65046 => x"ffffff",
   65047 => x"ffffff",
   65048 => x"ffffff",
   65049 => x"ffffff",
   65050 => x"ffffff",
   65051 => x"ffffff",
   65052 => x"ffffff",
   65053 => x"ffffff",
   65054 => x"ffffff",
   65055 => x"ffffff",
   65056 => x"ffffff",
   65057 => x"ffffff",
   65058 => x"ffffff",
   65059 => x"ffffff",
   65060 => x"ffffff",
   65061 => x"ffffff",
   65062 => x"ffffff",
   65063 => x"ffffff",
   65064 => x"ffffff",
   65065 => x"ffffff",
   65066 => x"ffffff",
   65067 => x"ffffff",
   65068 => x"ffffff",
   65069 => x"ffffff",
   65070 => x"ffffff",
   65071 => x"ffffff",
   65072 => x"ffffff",
   65073 => x"ffffff",
   65074 => x"ffffff",
   65075 => x"ffffff",
   65076 => x"ffffff",
   65077 => x"ffffff",
   65078 => x"ffffff",
   65079 => x"ffffff",
   65080 => x"ffffff",
   65081 => x"ffffff",
   65082 => x"ffffff",
   65083 => x"ffffff",
   65084 => x"ffffff",
   65085 => x"ffffff",
   65086 => x"ffffff",
   65087 => x"ffffff",
   65088 => x"ffffff",
   65089 => x"ffffff",
   65090 => x"ffffff",
   65091 => x"ffffff",
   65092 => x"ffffff",
   65093 => x"ffffff",
   65094 => x"ffffff",
   65095 => x"ffffff",
   65096 => x"ffffff",
   65097 => x"ffffff",
   65098 => x"ffffff",
   65099 => x"ffffff",
   65100 => x"ffffff",
   65101 => x"ffffff",
   65102 => x"ffffff",
   65103 => x"ffffff",
   65104 => x"ffffff",
   65105 => x"ffffff",
   65106 => x"ffffff",
   65107 => x"ffffff",
   65108 => x"ffffff",
   65109 => x"ffffff",
   65110 => x"ffffff",
   65111 => x"ffffff",
   65112 => x"ffffff",
   65113 => x"ffffff",
   65114 => x"ffffff",
   65115 => x"ffffff",
   65116 => x"ffffff",
   65117 => x"ffffff",
   65118 => x"ffffff",
   65119 => x"ffffff",
   65120 => x"ffffff",
   65121 => x"ffffff",
   65122 => x"ffffff",
   65123 => x"ffffff",
   65124 => x"ffffff",
   65125 => x"ffffff",
   65126 => x"ffffff",
   65127 => x"ffffff",
   65128 => x"ffffff",
   65129 => x"ffffff",
   65130 => x"ffffff",
   65131 => x"ffffff",
   65132 => x"ffffff",
   65133 => x"ffffff",
   65134 => x"ffffff",
   65135 => x"ffffff",
   65136 => x"ffffff",
   65137 => x"ffffff",
   65138 => x"ffffff",
   65139 => x"ffffff",
   65140 => x"ffffff",
   65141 => x"ffffff",
   65142 => x"ffffff",
   65143 => x"ffffff",
   65144 => x"ffffff",
   65145 => x"ffffff",
   65146 => x"ffffff",
   65147 => x"ffffff",
   65148 => x"ffffff",
   65149 => x"ffffff",
   65150 => x"ffffff",
   65151 => x"ffffff",
   65152 => x"ffffff",
   65153 => x"ffffff",
   65154 => x"ffffff",
   65155 => x"ffffff",
   65156 => x"ffffff",
   65157 => x"ffffff",
   65158 => x"ffffff",
   65159 => x"ffffff",
   65160 => x"ffffff",
   65161 => x"ffffff",
   65162 => x"ffffff",
   65163 => x"ffffff",
   65164 => x"ffffff",
   65165 => x"ffffff",
   65166 => x"ffffff",
   65167 => x"ffffff",
   65168 => x"ffffff",
   65169 => x"ffffff",
   65170 => x"ffffff",
   65171 => x"ffffff",
   65172 => x"ffffff",
   65173 => x"ffffff",
   65174 => x"ffffff",
   65175 => x"ffffff",
   65176 => x"ffffff",
   65177 => x"ffffff",
   65178 => x"ffffff",
   65179 => x"ffffff",
   65180 => x"ffffff",
   65181 => x"ffffff",
   65182 => x"ffffff",
   65183 => x"ffffff",
   65184 => x"ffffff",
   65185 => x"ffffff",
   65186 => x"ffffff",
   65187 => x"ffffff",
   65188 => x"ffffff",
   65189 => x"ffffff",
   65190 => x"ffffff",
   65191 => x"ffffff",
   65192 => x"ffffff",
   65193 => x"ffffff",
   65194 => x"ffffff",
   65195 => x"ffffff",
   65196 => x"ffffff",
   65197 => x"ffffff",
   65198 => x"ffffff",
   65199 => x"ffffff",
   65200 => x"ffffff",
   65201 => x"ffffff",
   65202 => x"ffffff",
   65203 => x"ffffff",
   65204 => x"ffffff",
   65205 => x"ffffff",
   65206 => x"ffffff",
   65207 => x"ffffff",
   65208 => x"ffffff",
   65209 => x"ffffff",
   65210 => x"ffffff",
   65211 => x"ffffff",
   65212 => x"ffffff",
   65213 => x"ffffff",
   65214 => x"ffffff",
   65215 => x"ffffff",
   65216 => x"ffffff",
   65217 => x"ffffff",
   65218 => x"ffffff",
   65219 => x"ffffff",
   65220 => x"ffffff",
   65221 => x"ffffff",
   65222 => x"ffffff",
   65223 => x"ffffff",
   65224 => x"ffffff",
   65225 => x"ffffff",
   65226 => x"ffffff",
   65227 => x"ffffff",
   65228 => x"ffffff",
   65229 => x"ffffff",
   65230 => x"ffffff",
   65231 => x"ffffff",
   65232 => x"ffffff",
   65233 => x"ffffff",
   65234 => x"ffffff",
   65235 => x"ffffff",
   65236 => x"ffffff",
   65237 => x"ffffff",
   65238 => x"ffffff",
   65239 => x"ffffff",
   65240 => x"ffffff",
   65241 => x"ffffff",
   65242 => x"ffffff",
   65243 => x"ffffff",
   65244 => x"ffffff",
   65245 => x"ffffff",
   65246 => x"ffffff",
   65247 => x"ffffff",
   65248 => x"ffffff",
   65249 => x"ffffff",
   65250 => x"ffffff",
   65251 => x"ffffff",
   65252 => x"ffffff",
   65253 => x"ffffff",
   65254 => x"ffffff",
   65255 => x"ffffff",
   65256 => x"ffffff",
   65257 => x"ffffff",
   65258 => x"ffffff",
   65259 => x"ffffff",
   65260 => x"ffffff",
   65261 => x"ffffff",
   65262 => x"ffffff",
   65263 => x"ffffff",
   65264 => x"ffffff",
   65265 => x"ffffff",
   65266 => x"ffffff",
   65267 => x"ffffff",
   65268 => x"ffffff",
   65269 => x"ffffff",
   65270 => x"ffffff",
   65271 => x"ffffff",
   65272 => x"ffffff",
   65273 => x"ffffff",
   65274 => x"ffffff",
   65275 => x"ffffff",
   65276 => x"ffffff",
   65277 => x"ffffff",
   65278 => x"ffffff",
   65279 => x"ffffff",
   65280 => x"ffffff",
   65281 => x"ffffff",
   65282 => x"ffffff",
   65283 => x"ffffff",
   65284 => x"ffffff",
   65285 => x"ffffff",
   65286 => x"ffffff",
   65287 => x"ffffff",
   65288 => x"ffffff",
   65289 => x"ffffff",
   65290 => x"ffffff",
   65291 => x"ffffff",
   65292 => x"ffffff",
   65293 => x"ffffff",
   65294 => x"ffffff",
   65295 => x"ffffff",
   65296 => x"ffffff",
   65297 => x"ffffff",
   65298 => x"ffffff",
   65299 => x"ffffff",
   65300 => x"ffffff",
   65301 => x"ffffff",
   65302 => x"ffffff",
   65303 => x"ffffff",
   65304 => x"ffffff",
   65305 => x"ffffff",
   65306 => x"ffffff",
   65307 => x"ffffff",
   65308 => x"ffffff",
   65309 => x"ffffff",
   65310 => x"ffffff",
   65311 => x"ffffff",
   65312 => x"ffffff",
   65313 => x"ffffff",
   65314 => x"ffffff",
   65315 => x"ffffff",
   65316 => x"ffffff",
   65317 => x"ffffff",
   65318 => x"ffffff",
   65319 => x"ffffff",
   65320 => x"ffffff",
   65321 => x"ffffff",
   65322 => x"ffffff",
   65323 => x"ffffff",
   65324 => x"ffffff",
   65325 => x"ffffff",
   65326 => x"ffffff",
   65327 => x"ffffff",
   65328 => x"ffffff",
   65329 => x"ffffff",
   65330 => x"ffffff",
   65331 => x"ffffff",
   65332 => x"ffffff",
   65333 => x"ffffff",
   65334 => x"ffffff",
   65335 => x"ffffff",
   65336 => x"ffffff",
   65337 => x"ffffff",
   65338 => x"ffffff",
   65339 => x"ffffff",
   65340 => x"ffffff",
   65341 => x"ffffff",
   65342 => x"ffffff",
   65343 => x"ffffff",
   65344 => x"ffffff",
   65345 => x"ffffff",
   65346 => x"ffffff",
   65347 => x"ffffff",
   65348 => x"ffffff",
   65349 => x"ffffff",
   65350 => x"ffffff",
   65351 => x"ffffff",
   65352 => x"ffffff",
   65353 => x"ffffff",
   65354 => x"ffffff",
   65355 => x"ffffff",
   65356 => x"ffffff",
   65357 => x"ffffff",
   65358 => x"ffffff",
   65359 => x"ffffff",
   65360 => x"ffffff",
   65361 => x"ffffff",
   65362 => x"ffffff",
   65363 => x"ffffff",
   65364 => x"ffffff",
   65365 => x"ffffff",
   65366 => x"ffffff",
   65367 => x"ffffff",
   65368 => x"ffffff",
   65369 => x"ffffff",
   65370 => x"ffffff",
   65371 => x"ffffff",
   65372 => x"ffffff",
   65373 => x"ffffff",
   65374 => x"ffffff",
   65375 => x"ffffff",
   65376 => x"ffffff",
   65377 => x"ffffff",
   65378 => x"ffffff",
   65379 => x"ffffff",
   65380 => x"ffffff",
   65381 => x"ffffff",
   65382 => x"ffffff",
   65383 => x"ffffff",
   65384 => x"ffffff",
   65385 => x"ffffff",
   65386 => x"ffffff",
   65387 => x"ffffff",
   65388 => x"ffffff",
   65389 => x"ffffff",
   65390 => x"ffffff",
   65391 => x"ffffff",
   65392 => x"ffffff",
   65393 => x"ffffff",
   65394 => x"ffffff",
   65395 => x"ffffff",
   65396 => x"ffffff",
   65397 => x"ffffff",
   65398 => x"ffffff",
   65399 => x"ffffff",
   65400 => x"ffffff",
   65401 => x"ffffff",
   65402 => x"ffffff",
   65403 => x"ffffff",
   65404 => x"ffffff",
   65405 => x"ffffff",
   65406 => x"ffffff",
   65407 => x"ffffff",
   65408 => x"ffffff",
   65409 => x"ffffff",
   65410 => x"ffffff",
   65411 => x"ffffff",
   65412 => x"ffffff",
   65413 => x"ffffff",
   65414 => x"ffffff",
   65415 => x"ffffff",
   65416 => x"ffffff",
   65417 => x"ffffff",
   65418 => x"ffffff",
   65419 => x"ffffff",
   65420 => x"ffffff",
   65421 => x"ffffff",
   65422 => x"ffffff",
   65423 => x"ffffff",
   65424 => x"ffffff",
   65425 => x"ffffff",
   65426 => x"ffffff",
   65427 => x"ffffff",
   65428 => x"ffffff",
   65429 => x"ffffff",
   65430 => x"ffffff",
   65431 => x"ffffff",
   65432 => x"ffffff",
   65433 => x"ffffff",
   65434 => x"ffffff",
   65435 => x"ffffff",
   65436 => x"ffffff",
   65437 => x"ffffff",
   65438 => x"ffffff",
   65439 => x"ffffff",
   65440 => x"ffffff",
   65441 => x"ffffff",
   65442 => x"ffffff",
   65443 => x"ffffff",
   65444 => x"ffffff",
   65445 => x"ffffff",
   65446 => x"ffffff",
   65447 => x"ffffff",
   65448 => x"ffffff",
   65449 => x"ffffff",
   65450 => x"ffffff",
   65451 => x"ffffff",
   65452 => x"ffffff",
   65453 => x"ffffff",
   65454 => x"ffffff",
   65455 => x"ffffff",
   65456 => x"ffffff",
   65457 => x"ffffff",
   65458 => x"ffffff",
   65459 => x"ffffff",
   65460 => x"ffffff",
   65461 => x"ffffff",
   65462 => x"ffffff",
   65463 => x"ffffff",
   65464 => x"ffffff",
   65465 => x"ffffff",
   65466 => x"ffffff",
   65467 => x"ffffff",
   65468 => x"ffffff",
   65469 => x"ffffff",
   65470 => x"ffffff",
   65471 => x"ffffff",
   65472 => x"ffffff",
   65473 => x"ffffff",
   65474 => x"ffffff",
   65475 => x"ffffff",
   65476 => x"ffffff",
   65477 => x"ffffff",
   65478 => x"ffffff",
   65479 => x"ffffff",
   65480 => x"ffffff",
   65481 => x"ffffff",
   65482 => x"ffffff",
   65483 => x"ffffff",
   65484 => x"ffffff",
   65485 => x"ffffff",
   65486 => x"ffffff",
   65487 => x"ffffff",
   65488 => x"ffffff",
   65489 => x"ffffff",
   65490 => x"ffffff",
   65491 => x"ffffff",
   65492 => x"ffffff",
   65493 => x"ffffff",
   65494 => x"ffffff",
   65495 => x"ffffff",
   65496 => x"ffffff",
   65497 => x"ffffff",
   65498 => x"ffffff",
   65499 => x"ffffff",
   65500 => x"ffffff",
   65501 => x"ffffff",
   65502 => x"ffffff",
   65503 => x"ffffff",
   65504 => x"ffffff",
   65505 => x"ffffff",
   65506 => x"ffffff",
   65507 => x"ffffff",
   65508 => x"ffffff",
   65509 => x"ffffff",
   65510 => x"ffffff",
   65511 => x"ffffff",
   65512 => x"ffffff",
   65513 => x"ffffff",
   65514 => x"ffffff",
   65515 => x"ffffff",
   65516 => x"ffffff",
   65517 => x"ffffff",
   65518 => x"ffffff",
   65519 => x"ffffff",
   65520 => x"ffffff",
   65521 => x"ffffff",
   65522 => x"ffffff",
   65523 => x"ffffff",
   65524 => x"ffffff",
   65525 => x"ffffff",
   65526 => x"ffffff",
   65527 => x"ffffff",
   65528 => x"ffffff",
   65529 => x"ffffff",
   65530 => x"ffffff",
   65531 => x"ffffff",
   65532 => x"ffffff",
   65533 => x"ffffff",
   65534 => x"ffffff",
   65535 => x"ffffff",
   65536 => x"ffffff",
   65537 => x"ffffff",
   65538 => x"ffffff",
   65539 => x"ffffff",
   65540 => x"ffffff",
   65541 => x"ffffff",
   65542 => x"ffffff",
   65543 => x"ffffff",
   65544 => x"ffffff",
   65545 => x"ffffff",
   65546 => x"ffffff",
   65547 => x"ffffff",
   65548 => x"ffffff",
   65549 => x"ffffff",
   65550 => x"ffffff",
   65551 => x"ffffff",
   65552 => x"ffffff",
   65553 => x"ffffff",
   65554 => x"ffffff",
   65555 => x"ffffff",
   65556 => x"ffffff",
   65557 => x"ffffff",
   65558 => x"ffffff",
   65559 => x"ffffff",
   65560 => x"ffffff",
   65561 => x"ffffff",
   65562 => x"ffffff",
   65563 => x"ffffff",
   65564 => x"ffffff",
   65565 => x"ffffff",
   65566 => x"ffffff",
   65567 => x"ffffff",
   65568 => x"ffffff",
   65569 => x"ffffff",
   65570 => x"ffffff",
   65571 => x"ffffff",
   65572 => x"ffffff",
   65573 => x"ffffff",
   65574 => x"ffffff",
   65575 => x"ffffff",
   65576 => x"ffffff",
   65577 => x"ffffff",
   65578 => x"ffffff",
   65579 => x"ffffff",
   65580 => x"ffffff",
   65581 => x"ffffff",
   65582 => x"ffffff",
   65583 => x"ffffff",
   65584 => x"ffffff",
   65585 => x"ffffff",
   65586 => x"ffffff",
   65587 => x"ffffff",
   65588 => x"ffffff",
   65589 => x"ffffff",
   65590 => x"ffffff",
   65591 => x"ffffff",
   65592 => x"ffffff",
   65593 => x"ffffff",
   65594 => x"ffffff",
   65595 => x"ffffff",
   65596 => x"ffffff",
   65597 => x"ffffff",
   65598 => x"ffffff",
   65599 => x"ffffff",
   65600 => x"ffffff",
   65601 => x"ffffff",
   65602 => x"ffffff",
   65603 => x"ffffff",
   65604 => x"ffffff",
   65605 => x"ffffff",
   65606 => x"ffffff",
   65607 => x"ffffff",
   65608 => x"ffffff",
   65609 => x"ffffff",
   65610 => x"ffffff",
   65611 => x"ffffff",
   65612 => x"ffffff",
   65613 => x"ffffff",
   65614 => x"ffffff",
   65615 => x"ffffff",
   65616 => x"ffffff",
   65617 => x"ffffff",
   65618 => x"ffffff",
   65619 => x"ffffff",
   65620 => x"ffffff",
   65621 => x"ffffff",
   65622 => x"ffffff",
   65623 => x"ffffff",
   65624 => x"ffffff",
   65625 => x"ffffff",
   65626 => x"ffffff",
   65627 => x"ffffff",
   65628 => x"ffffff",
   65629 => x"ffffff",
   65630 => x"ffffff",
   65631 => x"ffffff",
   65632 => x"ffffff",
   65633 => x"ffffff",
   65634 => x"ffffff",
   65635 => x"ffffff",
   65636 => x"ffffff",
   65637 => x"ffffff",
   65638 => x"ffffff",
   65639 => x"ffffff",
   65640 => x"ffffff",
   65641 => x"ffffff",
   65642 => x"ffffff",
   65643 => x"ffffff",
   65644 => x"ffffff",
   65645 => x"ffffff",
   65646 => x"ffffff",
   65647 => x"ffffff",
   65648 => x"ffffff",
   65649 => x"ffffff",
   65650 => x"ffffff",
   65651 => x"ffffff",
   65652 => x"ffffff",
   65653 => x"ffffff",
   65654 => x"ffffff",
   65655 => x"ffffff",
   65656 => x"ffffff",
   65657 => x"ffffff",
   65658 => x"ffffff",
   65659 => x"ffffff",
   65660 => x"ffffff",
   65661 => x"ffffff",
   65662 => x"ffffff",
   65663 => x"ffffff",
   65664 => x"ffffff",
   65665 => x"ffffff",
   65666 => x"ffffff",
   65667 => x"ffffff",
   65668 => x"ffffff",
   65669 => x"ffffff",
   65670 => x"ffffff",
   65671 => x"ffffff",
   65672 => x"ffffff",
   65673 => x"ffffff",
   65674 => x"ffffff",
   65675 => x"ffffff",
   65676 => x"ffffff",
   65677 => x"ffffff",
   65678 => x"ffffff",
   65679 => x"ffffff",
   65680 => x"ffffff",
   65681 => x"ffffff",
   65682 => x"ffffff",
   65683 => x"ffffff",
   65684 => x"ffffff",
   65685 => x"ffffff",
   65686 => x"ffffff",
   65687 => x"ffffff",
   65688 => x"ffffff",
   65689 => x"ffffff",
   65690 => x"ffffff",
   65691 => x"ffffff",
   65692 => x"ffffff",
   65693 => x"ffffff",
   65694 => x"ffffff",
   65695 => x"ffffff",
   65696 => x"ffffff",
   65697 => x"ffffff",
   65698 => x"ffffff",
   65699 => x"ffffff",
   65700 => x"ffffff",
   65701 => x"ffffff",
   65702 => x"ffffff",
   65703 => x"ffffff",
   65704 => x"ffffff",
   65705 => x"ffffff",
   65706 => x"ffffff",
   65707 => x"ffffff",
   65708 => x"ffffff",
   65709 => x"ffffff",
   65710 => x"ffffff",
   65711 => x"ffffff",
   65712 => x"ffffff",
   65713 => x"ffffff",
   65714 => x"ffffff",
   65715 => x"ffffff",
   65716 => x"ffffff",
   65717 => x"ffffff",
   65718 => x"ffffff",
   65719 => x"ffffff",
   65720 => x"ffffff",
   65721 => x"ffffff",
   65722 => x"ffffff",
   65723 => x"ffffff",
   65724 => x"ffffff",
   65725 => x"ffffff",
   65726 => x"ffffff",
   65727 => x"ffffff",
   65728 => x"ffffff",
   65729 => x"ffffff",
   65730 => x"ffffff",
   65731 => x"ffffff",
   65732 => x"ffffff",
   65733 => x"ffffff",
   65734 => x"ffffff",
   65735 => x"ffffff",
   65736 => x"ffffff",
   65737 => x"ffffff",
   65738 => x"ffffff",
   65739 => x"ffffff",
   65740 => x"ffffff",
   65741 => x"ffffff",
   65742 => x"ffffff",
   65743 => x"ffffff",
   65744 => x"ffffff",
   65745 => x"ffffff",
   65746 => x"ffffff",
   65747 => x"ffffff",
   65748 => x"ffffff",
   65749 => x"ffffff",
   65750 => x"ffffff",
   65751 => x"ffffff",
   65752 => x"ffffff",
   65753 => x"ffffff",
   65754 => x"ffffff",
   65755 => x"ffffff",
   65756 => x"ffffff",
   65757 => x"ffffff",
   65758 => x"ffffff",
   65759 => x"ffffff",
   65760 => x"ffffff",
   65761 => x"ffffff",
   65762 => x"ffffff",
   65763 => x"ffffff",
   65764 => x"ffffff",
   65765 => x"ffffff",
   65766 => x"ffffff",
   65767 => x"ffffff",
   65768 => x"ffffff",
   65769 => x"ffffff",
   65770 => x"ffffff",
   65771 => x"ffffff",
   65772 => x"ffffff",
   65773 => x"ffffff",
   65774 => x"ffffff",
   65775 => x"ffffff",
   65776 => x"ffffff",
   65777 => x"ffffff",
   65778 => x"ffffff",
   65779 => x"ffffff",
   65780 => x"ffffff",
   65781 => x"ffffff",
   65782 => x"ffffff",
   65783 => x"ffffff",
   65784 => x"ffffff",
   65785 => x"ffffff",
   65786 => x"ffffff",
   65787 => x"ffffff",
   65788 => x"ffffff",
   65789 => x"ffffff",
   65790 => x"ffffff",
   65791 => x"ffffff",
   65792 => x"ffffff",
   65793 => x"ffffff",
   65794 => x"ffffff",
   65795 => x"ffffff",
   65796 => x"ffffff",
   65797 => x"ffffff",
   65798 => x"ffffff",
   65799 => x"ffffff",
   65800 => x"ffffff",
   65801 => x"ffffff",
   65802 => x"ffffff",
   65803 => x"ffffff",
   65804 => x"ffffff",
   65805 => x"ffffff",
   65806 => x"ffffff",
   65807 => x"ffffff",
   65808 => x"ffffff",
   65809 => x"ffffff",
   65810 => x"ffffff",
   65811 => x"ffffff",
   65812 => x"ffffff",
   65813 => x"ffffff",
   65814 => x"ffffff",
   65815 => x"ffffff",
   65816 => x"ffffff",
   65817 => x"ffffff",
   65818 => x"ffffff",
   65819 => x"ffffff",
   65820 => x"ffffff",
   65821 => x"ffffff",
   65822 => x"ffffff",
   65823 => x"ffffff",
   65824 => x"ffffff",
   65825 => x"ffffff",
   65826 => x"ffffff",
   65827 => x"ffffff",
   65828 => x"ffffff",
   65829 => x"ffffff",
   65830 => x"ffffff",
   65831 => x"ffffff",
   65832 => x"ffffff",
   65833 => x"ffffff",
   65834 => x"ffffff",
   65835 => x"ffffff",
   65836 => x"ffffff",
   65837 => x"ffffff",
   65838 => x"ffffff",
   65839 => x"ffffff",
   65840 => x"ffffff",
   65841 => x"ffffff",
   65842 => x"ffffff",
   65843 => x"ffffff",
   65844 => x"ffffff",
   65845 => x"ffffff",
   65846 => x"ffffff",
   65847 => x"ffffff",
   65848 => x"ffffff",
   65849 => x"ffffff",
   65850 => x"ffffff",
   65851 => x"ffffff",
   65852 => x"ffffff",
   65853 => x"ffffff",
   65854 => x"ffffff",
   65855 => x"ffffff",
   65856 => x"ffffff",
   65857 => x"ffffff",
   65858 => x"ffffff",
   65859 => x"ffffff",
   65860 => x"ffffff",
   65861 => x"ffffff",
   65862 => x"ffffff",
   65863 => x"ffffff",
   65864 => x"ffffff",
   65865 => x"ffffff",
   65866 => x"ffffff",
   65867 => x"ffffff",
   65868 => x"ffffff",
   65869 => x"ffffff",
   65870 => x"ffffff",
   65871 => x"ffffff",
   65872 => x"ffffff",
   65873 => x"ffffff",
   65874 => x"ffffff",
   65875 => x"ffffff",
   65876 => x"ffffff",
   65877 => x"ffffff",
   65878 => x"ffffff",
   65879 => x"ffffff",
   65880 => x"ffffff",
   65881 => x"ffffff",
   65882 => x"ffffff",
   65883 => x"ffffff",
   65884 => x"ffffff",
   65885 => x"ffffff",
   65886 => x"ffffff",
   65887 => x"ffffff",
   65888 => x"ffffff",
   65889 => x"ffffff",
   65890 => x"ffffff",
   65891 => x"ffffff",
   65892 => x"ffffff",
   65893 => x"ffffff",
   65894 => x"ffffff",
   65895 => x"ffffff",
   65896 => x"ffffff",
   65897 => x"ffffff",
   65898 => x"ffffff",
   65899 => x"ffffff",
   65900 => x"ffffff",
   65901 => x"ffffff",
   65902 => x"ffffff",
   65903 => x"ffffff",
   65904 => x"ffffff",
   65905 => x"ffffff",
   65906 => x"ffffff",
   65907 => x"ffffff",
   65908 => x"ffffff",
   65909 => x"ffffff",
   65910 => x"ffffff",
   65911 => x"ffffff",
   65912 => x"ffffff",
   65913 => x"ffffff",
   65914 => x"ffffff",
   65915 => x"ffffff",
   65916 => x"ffffff",
   65917 => x"ffffff",
   65918 => x"ffffff",
   65919 => x"ffffff",
   65920 => x"ffffff",
   65921 => x"ffffff",
   65922 => x"ffffff",
   65923 => x"ffffff",
   65924 => x"ffffff",
   65925 => x"ffffff",
   65926 => x"ffffff",
   65927 => x"ffffff",
   65928 => x"ffffff",
   65929 => x"ffffff",
   65930 => x"ffffff",
   65931 => x"ffffff",
   65932 => x"ffffff",
   65933 => x"ffffff",
   65934 => x"ffffff",
   65935 => x"ffffff",
   65936 => x"ffffff",
   65937 => x"ffffff",
   65938 => x"ffffff",
   65939 => x"ffffff",
   65940 => x"ffffff",
   65941 => x"ffffff",
   65942 => x"ffffff",
   65943 => x"ffffff",
   65944 => x"ffffff",
   65945 => x"ffffff",
   65946 => x"ffffff",
   65947 => x"ffffff",
   65948 => x"ffffff",
   65949 => x"ffffff",
   65950 => x"ffffff",
   65951 => x"ffffff",
   65952 => x"ffffff",
   65953 => x"ffffff",
   65954 => x"ffffff",
   65955 => x"ffffff",
   65956 => x"ffffff",
   65957 => x"ffffff",
   65958 => x"ffffff",
   65959 => x"ffffff",
   65960 => x"ffffff",
   65961 => x"ffffff",
   65962 => x"ffffff",
   65963 => x"ffffff",
   65964 => x"ffffff",
   65965 => x"ffffff",
   65966 => x"ffffff",
   65967 => x"ffffff",
   65968 => x"ffffff",
   65969 => x"ffffff",
   65970 => x"ffffff",
   65971 => x"ffffff",
   65972 => x"ffffff",
   65973 => x"ffffff",
   65974 => x"ffffff",
   65975 => x"ffffff",
   65976 => x"ffffff",
   65977 => x"ffffff",
   65978 => x"ffffff",
   65979 => x"ffffff",
   65980 => x"ffffff",
   65981 => x"ffffff",
   65982 => x"ffffff",
   65983 => x"ffffff",
   65984 => x"ffffff",
   65985 => x"ffffff",
   65986 => x"ffffff",
   65987 => x"ffffff",
   65988 => x"ffffff",
   65989 => x"ffffff",
   65990 => x"ffffff",
   65991 => x"ffffff",
   65992 => x"ffffff",
   65993 => x"ffffff",
   65994 => x"ffffff",
   65995 => x"ffffff",
   65996 => x"ffffff",
   65997 => x"ffffff",
   65998 => x"ffffff",
   65999 => x"ffffff",
   66000 => x"ffffff",
   66001 => x"ffffff",
   66002 => x"ffffff",
   66003 => x"ffffff",
   66004 => x"ffffff",
   66005 => x"ffffff",
   66006 => x"ffffff",
   66007 => x"ffffff",
   66008 => x"ffffff",
   66009 => x"ffffff",
   66010 => x"ffffff",
   66011 => x"ffffff",
   66012 => x"ffffff",
   66013 => x"ffffff",
   66014 => x"ffffff",
   66015 => x"ffffff",
   66016 => x"ffffff",
   66017 => x"ffffff",
   66018 => x"ffffff",
   66019 => x"ffffff",
   66020 => x"ffffff",
   66021 => x"ffffff",
   66022 => x"ffffff",
   66023 => x"ffffff",
   66024 => x"ffffff",
   66025 => x"ffffff",
   66026 => x"ffffff",
   66027 => x"ffffff",
   66028 => x"ffffff",
   66029 => x"ffffff",
   66030 => x"ffffff",
   66031 => x"ffffff",
   66032 => x"ffffff",
   66033 => x"ffffff",
   66034 => x"ffffff",
   66035 => x"ffffff",
   66036 => x"ffffff",
   66037 => x"ffffff",
   66038 => x"ffffff",
   66039 => x"ffffff",
   66040 => x"ffffff",
   66041 => x"ffffff",
   66042 => x"ffffff",
   66043 => x"ffffff",
   66044 => x"ffffff",
   66045 => x"ffffff",
   66046 => x"ffffff",
   66047 => x"ffffff",
   66048 => x"ffffff",
   66049 => x"ffffff",
   66050 => x"ffffff",
   66051 => x"ffffff",
   66052 => x"ffffff",
   66053 => x"ffffff",
   66054 => x"ffffff",
   66055 => x"ffffff",
   66056 => x"ffffff",
   66057 => x"ffffff",
   66058 => x"ffffff",
   66059 => x"ffffff",
   66060 => x"ffffff",
   66061 => x"ffffff",
   66062 => x"ffffff",
   66063 => x"ffffff",
   66064 => x"ffffff",
   66065 => x"ffffff",
   66066 => x"ffffff",
   66067 => x"ffffff",
   66068 => x"ffffff",
   66069 => x"ffffff",
   66070 => x"ffffff",
   66071 => x"ffffff",
   66072 => x"ffffff",
   66073 => x"ffffff",
   66074 => x"ffffff",
   66075 => x"ffffff",
   66076 => x"ffffff",
   66077 => x"ffffff",
   66078 => x"ffffff",
   66079 => x"ffffff",
   66080 => x"ffffff",
   66081 => x"ffffff",
   66082 => x"ffffff",
   66083 => x"ffffff",
   66084 => x"ffffff",
   66085 => x"ffffff",
   66086 => x"ffffff",
   66087 => x"ffffff",
   66088 => x"ffffff",
   66089 => x"ffffff",
   66090 => x"ffffff",
   66091 => x"ffffff",
   66092 => x"ffffff",
   66093 => x"ffffff",
   66094 => x"ffffff",
   66095 => x"ffffff",
   66096 => x"ffffff",
   66097 => x"ffffff",
   66098 => x"ffffff",
   66099 => x"ffffff",
   66100 => x"ffffff",
   66101 => x"ffffff",
   66102 => x"ffffff",
   66103 => x"ffffff",
   66104 => x"ffffff",
   66105 => x"ffffff",
   66106 => x"ffffff",
   66107 => x"ffffff",
   66108 => x"ffffff",
   66109 => x"ffffff",
   66110 => x"ffffff",
   66111 => x"ffffff",
   66112 => x"ffffff",
   66113 => x"ffffff",
   66114 => x"ffffff",
   66115 => x"ffffff",
   66116 => x"ffffff",
   66117 => x"ffffff",
   66118 => x"ffffff",
   66119 => x"ffffff",
   66120 => x"ffffff",
   66121 => x"ffffff",
   66122 => x"ffffff",
   66123 => x"ffffff",
   66124 => x"ffffff",
   66125 => x"ffffff",
   66126 => x"ffffff",
   66127 => x"ffffff",
   66128 => x"ffffff",
   66129 => x"ffffff",
   66130 => x"ffffff",
   66131 => x"ffffff",
   66132 => x"ffffff",
   66133 => x"ffffff",
   66134 => x"ffffff",
   66135 => x"ffffff",
   66136 => x"ffffff",
   66137 => x"ffffff",
   66138 => x"ffffff",
   66139 => x"ffffff",
   66140 => x"ffffff",
   66141 => x"ffffff",
   66142 => x"ffffff",
   66143 => x"ffffff",
   66144 => x"ffffff",
   66145 => x"ffffff",
   66146 => x"ffffff",
   66147 => x"ffffff",
   66148 => x"ffffff",
   66149 => x"ffffff",
   66150 => x"ffffff",
   66151 => x"ffffff",
   66152 => x"ffffff",
   66153 => x"ffffff",
   66154 => x"ffffff",
   66155 => x"ffffff",
   66156 => x"ffffff",
   66157 => x"ffffff",
   66158 => x"ffffff",
   66159 => x"ffffff",
   66160 => x"ffffff",
   66161 => x"ffffff",
   66162 => x"ffffff",
   66163 => x"ffffff",
   66164 => x"ffffff",
   66165 => x"ffffff",
   66166 => x"ffffff",
   66167 => x"ffffff",
   66168 => x"ffffff",
   66169 => x"ffffff",
   66170 => x"ffffff",
   66171 => x"ffffff",
   66172 => x"ffffff",
   66173 => x"ffffff",
   66174 => x"ffffff",
   66175 => x"ffffff",
   66176 => x"ffffff",
   66177 => x"ffffff",
   66178 => x"ffffff",
   66179 => x"ffffff",
   66180 => x"ffffff",
   66181 => x"ffffff",
   66182 => x"ffffff",
   66183 => x"ffffff",
   66184 => x"ffffff",
   66185 => x"ffffff",
   66186 => x"ffffff",
   66187 => x"ffffff",
   66188 => x"ffffff",
   66189 => x"ffffff",
   66190 => x"ffffff",
   66191 => x"ffffff",
   66192 => x"ffffff",
   66193 => x"ffffff",
   66194 => x"ffffff",
   66195 => x"ffffff",
   66196 => x"ffffff",
   66197 => x"ffffff",
   66198 => x"ffffff",
   66199 => x"ffffff",
   66200 => x"ffffff",
   66201 => x"ffffff",
   66202 => x"ffffff",
   66203 => x"ffffff",
   66204 => x"ffffff",
   66205 => x"ffffff",
   66206 => x"ffffff",
   66207 => x"ffffff",
   66208 => x"ffffff",
   66209 => x"ffffff",
   66210 => x"ffffff",
   66211 => x"ffffff",
   66212 => x"ffffff",
   66213 => x"ffffff",
   66214 => x"ffffff",
   66215 => x"ffffff",
   66216 => x"ffffff",
   66217 => x"ffffff",
   66218 => x"ffffff",
   66219 => x"ffffff",
   66220 => x"ffffff",
   66221 => x"ffffff",
   66222 => x"ffffff",
   66223 => x"ffffff",
   66224 => x"ffffff",
   66225 => x"ffffff",
   66226 => x"ffffff",
   66227 => x"ffffff",
   66228 => x"ffffff",
   66229 => x"ffffff",
   66230 => x"ffffff",
   66231 => x"ffffff",
   66232 => x"ffffff",
   66233 => x"ffffff",
   66234 => x"ffffff",
   66235 => x"ffffff",
   66236 => x"ffffff",
   66237 => x"ffffff",
   66238 => x"ffffff",
   66239 => x"ffffff",
   66240 => x"ffffff",
   66241 => x"ffffff",
   66242 => x"ffffff",
   66243 => x"ffffff",
   66244 => x"ffffff",
   66245 => x"ffffff",
   66246 => x"ffffff",
   66247 => x"ffffff",
   66248 => x"ffffff",
   66249 => x"ffffff",
   66250 => x"ffffff",
   66251 => x"ffffff",
   66252 => x"ffffff",
   66253 => x"ffffff",
   66254 => x"ffffff",
   66255 => x"ffffff",
   66256 => x"ffffff",
   66257 => x"ffffff",
   66258 => x"ffffff",
   66259 => x"ffffff",
   66260 => x"ffffff",
   66261 => x"ffffff",
   66262 => x"ffffff",
   66263 => x"ffffff",
   66264 => x"ffffff",
   66265 => x"ffffff",
   66266 => x"ffffff",
   66267 => x"ffffff",
   66268 => x"ffffff",
   66269 => x"ffffff",
   66270 => x"ffffff",
   66271 => x"ffffff",
   66272 => x"ffffff",
   66273 => x"ffffff",
   66274 => x"ffffff",
   66275 => x"ffffff",
   66276 => x"ffffff",
   66277 => x"ffffff",
   66278 => x"ffffff",
   66279 => x"ffffff",
   66280 => x"ffffff",
   66281 => x"ffffff",
   66282 => x"ffffff",
   66283 => x"ffffff",
   66284 => x"ffffff",
   66285 => x"ffffff",
   66286 => x"ffffff",
   66287 => x"ffffff",
   66288 => x"ffffff",
   66289 => x"ffffff",
   66290 => x"ffffff",
   66291 => x"ffffff",
   66292 => x"ffffff",
   66293 => x"ffffff",
   66294 => x"ffffff",
   66295 => x"ffffff",
   66296 => x"ffffff",
   66297 => x"ffffff",
   66298 => x"ffffff",
   66299 => x"ffffff",
   66300 => x"ffffff",
   66301 => x"ffffff",
   66302 => x"ffffff",
   66303 => x"ffffff",
   66304 => x"ffffff",
   66305 => x"ffffff",
   66306 => x"ffffff",
   66307 => x"ffffff",
   66308 => x"ffffff",
   66309 => x"ffffff",
   66310 => x"ffffff",
   66311 => x"ffffff",
   66312 => x"ffffff",
   66313 => x"ffffff",
   66314 => x"ffffff",
   66315 => x"ffffff",
   66316 => x"ffffff",
   66317 => x"ffffff",
   66318 => x"ffffff",
   66319 => x"ffffff",
   66320 => x"ffffff",
   66321 => x"ffffff",
   66322 => x"ffffff",
   66323 => x"ffffff",
   66324 => x"ffffff",
   66325 => x"ffffff",
   66326 => x"ffffff",
   66327 => x"ffffff",
   66328 => x"ffffff",
   66329 => x"ffffff",
   66330 => x"ffffff",
   66331 => x"ffffff",
   66332 => x"ffffff",
   66333 => x"ffffff",
   66334 => x"ffffff",
   66335 => x"ffffff",
   66336 => x"ffffff",
   66337 => x"ffffff",
   66338 => x"ffffff",
   66339 => x"ffffff",
   66340 => x"ffffff",
   66341 => x"ffffff",
   66342 => x"ffffff",
   66343 => x"ffffff",
   66344 => x"ffffff",
   66345 => x"ffffff",
   66346 => x"ffffff",
   66347 => x"ffffff",
   66348 => x"ffffff",
   66349 => x"ffffff",
   66350 => x"ffffff",
   66351 => x"ffffff",
   66352 => x"ffffff",
   66353 => x"ffffff",
   66354 => x"ffffff",
   66355 => x"ffffff",
   66356 => x"ffffff",
   66357 => x"ffffff",
   66358 => x"ffffff",
   66359 => x"ffffff",
   66360 => x"ffffff",
   66361 => x"ffffff",
   66362 => x"ffffff",
   66363 => x"ffffff",
   66364 => x"ffffff",
   66365 => x"ffffff",
   66366 => x"ffffff",
   66367 => x"ffffff",
   66368 => x"ffffff",
   66369 => x"ffffff",
   66370 => x"ffffff",
   66371 => x"ffffff",
   66372 => x"ffffff",
   66373 => x"ffffff",
   66374 => x"ffffff",
   66375 => x"ffffff",
   66376 => x"ffffff",
   66377 => x"ffffff",
   66378 => x"ffffff",
   66379 => x"ffffff",
   66380 => x"ffffff",
   66381 => x"ffffff",
   66382 => x"ffffff",
   66383 => x"ffffff",
   66384 => x"ffffff",
   66385 => x"ffffff",
   66386 => x"ffffff",
   66387 => x"ffffff",
   66388 => x"ffffff",
   66389 => x"ffffff",
   66390 => x"ffffff",
   66391 => x"ffffff",
   66392 => x"ffffff",
   66393 => x"ffffff",
   66394 => x"ffffff",
   66395 => x"ffffff",
   66396 => x"ffffff",
   66397 => x"ffffff",
   66398 => x"ffffff",
   66399 => x"ffffff",
   66400 => x"ffffff",
   66401 => x"ffffff",
   66402 => x"ffffff",
   66403 => x"ffffff",
   66404 => x"ffffff",
   66405 => x"ffffff",
   66406 => x"ffffff",
   66407 => x"ffffff",
   66408 => x"ffffff",
   66409 => x"ffffff",
   66410 => x"ffffff",
   66411 => x"ffffff",
   66412 => x"ffffff",
   66413 => x"ffffff",
   66414 => x"ffffff",
   66415 => x"ffffff",
   66416 => x"ffffff",
   66417 => x"ffffff",
   66418 => x"ffffff",
   66419 => x"ffffff",
   66420 => x"ffffff",
   66421 => x"ffffff",
   66422 => x"ffffff",
   66423 => x"ffffff",
   66424 => x"ffffff",
   66425 => x"ffffff",
   66426 => x"ffffff",
   66427 => x"ffffff",
   66428 => x"ffffff",
   66429 => x"ffffff",
   66430 => x"ffffff",
   66431 => x"ffffff",
   66432 => x"ffffff",
   66433 => x"ffffff",
   66434 => x"ffffff",
   66435 => x"ffffff",
   66436 => x"ffffff",
   66437 => x"ffffff",
   66438 => x"ffffff",
   66439 => x"ffffff",
   66440 => x"ffffff",
   66441 => x"ffffff",
   66442 => x"ffffff",
   66443 => x"ffffff",
   66444 => x"ffffff",
   66445 => x"ffffff",
   66446 => x"ffffff",
   66447 => x"ffffff",
   66448 => x"ffffff",
   66449 => x"ffffff",
   66450 => x"ffffff",
   66451 => x"ffffff",
   66452 => x"ffffff",
   66453 => x"ffffff",
   66454 => x"ffffff",
   66455 => x"ffffff",
   66456 => x"ffffff",
   66457 => x"ffffff",
   66458 => x"ffffff",
   66459 => x"ffffff",
   66460 => x"ffffff",
   66461 => x"ffffff",
   66462 => x"ffffff",
   66463 => x"ffffff",
   66464 => x"ffffff",
   66465 => x"ffffff",
   66466 => x"ffffff",
   66467 => x"ffffff",
   66468 => x"ffffff",
   66469 => x"ffffff",
   66470 => x"ffffff",
   66471 => x"ffffff",
   66472 => x"ffffff",
   66473 => x"ffffff",
   66474 => x"ffffff",
   66475 => x"ffffff",
   66476 => x"ffffff",
   66477 => x"ffffff",
   66478 => x"ffffff",
   66479 => x"ffffff",
   66480 => x"ffffff",
   66481 => x"ffffff",
   66482 => x"ffffff",
   66483 => x"ffffff",
   66484 => x"ffffff",
   66485 => x"ffffff",
   66486 => x"ffffff",
   66487 => x"ffffff",
   66488 => x"ffffff",
   66489 => x"ffffff",
   66490 => x"ffffff",
   66491 => x"ffffff",
   66492 => x"ffffff",
   66493 => x"ffffff",
   66494 => x"ffffff",
   66495 => x"ffffff",
   66496 => x"ffffff",
   66497 => x"ffffff",
   66498 => x"ffffff",
   66499 => x"ffffff",
   66500 => x"ffffff",
   66501 => x"ffffff",
   66502 => x"ffffff",
   66503 => x"ffffff",
   66504 => x"ffffff",
   66505 => x"ffffff",
   66506 => x"ffffff",
   66507 => x"ffffff",
   66508 => x"ffffff",
   66509 => x"ffffff",
   66510 => x"ffffff",
   66511 => x"ffffff",
   66512 => x"ffffff",
   66513 => x"ffffff",
   66514 => x"ffffff",
   66515 => x"ffffff",
   66516 => x"ffffff",
   66517 => x"ffffff",
   66518 => x"ffffff",
   66519 => x"ffffff",
   66520 => x"ffffff",
   66521 => x"ffffff",
   66522 => x"ffffff",
   66523 => x"ffffff",
   66524 => x"ffffff",
   66525 => x"ffffff",
   66526 => x"ffffff",
   66527 => x"ffffff",
   66528 => x"ffffff",
   66529 => x"ffffff",
   66530 => x"ffffff",
   66531 => x"ffffff",
   66532 => x"ffffff",
   66533 => x"ffffff",
   66534 => x"ffffff",
   66535 => x"ffffff",
   66536 => x"ffffff",
   66537 => x"ffffff",
   66538 => x"ffffff",
   66539 => x"ffffff",
   66540 => x"ffffff",
   66541 => x"ffffff",
   66542 => x"ffffff",
   66543 => x"ffffff",
   66544 => x"ffffff",
   66545 => x"ffffff",
   66546 => x"ffffff",
   66547 => x"ffffff",
   66548 => x"ffffff",
   66549 => x"ffffff",
   66550 => x"ffffff",
   66551 => x"ffffff",
   66552 => x"ffffff",
   66553 => x"ffffff",
   66554 => x"ffffff",
   66555 => x"ffffff",
   66556 => x"ffffff",
   66557 => x"ffffff",
   66558 => x"ffffff",
   66559 => x"ffffff",
   66560 => x"ffffff",
   66561 => x"ffffff",
   66562 => x"ffffff",
   66563 => x"ffffff",
   66564 => x"ffffff",
   66565 => x"ffffff",
   66566 => x"ffffff",
   66567 => x"ffffff",
   66568 => x"ffffff",
   66569 => x"ffffff",
   66570 => x"ffffff",
   66571 => x"ffffff",
   66572 => x"ffffff",
   66573 => x"ffffff",
   66574 => x"ffffff",
   66575 => x"ffffff",
   66576 => x"ffffff",
   66577 => x"ffffff",
   66578 => x"ffffff",
   66579 => x"ffffff",
   66580 => x"ffffff",
   66581 => x"ffffff",
   66582 => x"ffffff",
   66583 => x"ffffff",
   66584 => x"ffffff",
   66585 => x"ffffff",
   66586 => x"ffffff",
   66587 => x"ffffff",
   66588 => x"ffffff",
   66589 => x"ffffff",
   66590 => x"ffffff",
   66591 => x"ffffff",
   66592 => x"ffffff",
   66593 => x"ffffff",
   66594 => x"ffffff",
   66595 => x"ffffff",
   66596 => x"ffffff",
   66597 => x"ffffff",
   66598 => x"ffffff",
   66599 => x"ffffff",
   66600 => x"ffffff",
   66601 => x"ffffff",
   66602 => x"ffffff",
   66603 => x"ffffff",
   66604 => x"ffffff",
   66605 => x"ffffff",
   66606 => x"ffffff",
   66607 => x"ffffff",
   66608 => x"ffffff",
   66609 => x"ffffff",
   66610 => x"ffffff",
   66611 => x"ffffff",
   66612 => x"ffffff",
   66613 => x"ffffff",
   66614 => x"ffffff",
   66615 => x"ffffff",
   66616 => x"ffffff",
   66617 => x"ffffff",
   66618 => x"ffffff",
   66619 => x"ffffff",
   66620 => x"ffffff",
   66621 => x"ffffff",
   66622 => x"ffffff",
   66623 => x"ffffff",
   66624 => x"ffffff",
   66625 => x"ffffff",
   66626 => x"ffffff",
   66627 => x"ffffff",
   66628 => x"ffffff",
   66629 => x"ffffff",
   66630 => x"ffffff",
   66631 => x"ffffff",
   66632 => x"ffffff",
   66633 => x"ffffff",
   66634 => x"ffffff",
   66635 => x"ffffff",
   66636 => x"ffffff",
   66637 => x"ffffff",
   66638 => x"ffffff",
   66639 => x"ffffff",
   66640 => x"ffffff",
   66641 => x"ffffff",
   66642 => x"ffffff",
   66643 => x"ffffff",
   66644 => x"ffffff",
   66645 => x"ffffff",
   66646 => x"ffffff",
   66647 => x"ffffff",
   66648 => x"ffffff",
   66649 => x"ffffff",
   66650 => x"ffffff",
   66651 => x"ffffff",
   66652 => x"ffffff",
   66653 => x"ffffff",
   66654 => x"ffffff",
   66655 => x"ffffff",
   66656 => x"ffffff",
   66657 => x"ffffff",
   66658 => x"ffffff",
   66659 => x"ffffff",
   66660 => x"ffffff",
   66661 => x"ffffff",
   66662 => x"ffffff",
   66663 => x"ffffff",
   66664 => x"ffffff",
   66665 => x"ffffff",
   66666 => x"ffffff",
   66667 => x"ffffff",
   66668 => x"ffffff",
   66669 => x"ffffff",
   66670 => x"ffffff",
   66671 => x"ffffff",
   66672 => x"ffffff",
   66673 => x"ffffff",
   66674 => x"ffffff",
   66675 => x"ffffff",
   66676 => x"ffffff",
   66677 => x"ffffff",
   66678 => x"ffffff",
   66679 => x"ffffff",
   66680 => x"ffffff",
   66681 => x"ffffff",
   66682 => x"ffffff",
   66683 => x"ffffff",
   66684 => x"ffffff",
   66685 => x"ffffff",
   66686 => x"ffffff",
   66687 => x"ffffff",
   66688 => x"ffffff",
   66689 => x"ffffff",
   66690 => x"ffffff",
   66691 => x"ffffff",
   66692 => x"ffffff",
   66693 => x"ffffff",
   66694 => x"ffffff",
   66695 => x"ffffff",
   66696 => x"ffffff",
   66697 => x"ffffff",
   66698 => x"ffffff",
   66699 => x"ffffff",
   66700 => x"ffffff",
   66701 => x"ffffff",
   66702 => x"ffffff",
   66703 => x"ffffff",
   66704 => x"ffffff",
   66705 => x"ffffff",
   66706 => x"ffffff",
   66707 => x"ffffff",
   66708 => x"ffffff",
   66709 => x"ffffff",
   66710 => x"ffffff",
   66711 => x"ffffff",
   66712 => x"ffffff",
   66713 => x"ffffff",
   66714 => x"ffffff",
   66715 => x"ffffff",
   66716 => x"ffffff",
   66717 => x"ffffff",
   66718 => x"ffffff",
   66719 => x"ffffff",
   66720 => x"ffffff",
   66721 => x"ffffff",
   66722 => x"ffffff",
   66723 => x"ffffff",
   66724 => x"ffffff",
   66725 => x"ffffff",
   66726 => x"ffffff",
   66727 => x"ffffff",
   66728 => x"ffffff",
   66729 => x"ffffff",
   66730 => x"ffffff",
   66731 => x"ffffff",
   66732 => x"ffffff",
   66733 => x"ffffff",
   66734 => x"ffffff",
   66735 => x"ffffff",
   66736 => x"ffffff",
   66737 => x"ffffff",
   66738 => x"ffffff",
   66739 => x"ffffff",
   66740 => x"ffffff",
   66741 => x"ffffff",
   66742 => x"ffffff",
   66743 => x"ffffff",
   66744 => x"ffffff",
   66745 => x"ffffff",
   66746 => x"ffffff",
   66747 => x"ffffff",
   66748 => x"ffffff",
   66749 => x"ffffff",
   66750 => x"ffffff",
   66751 => x"ffffff",
   66752 => x"ffffff",
   66753 => x"ffffff",
   66754 => x"ffffff",
   66755 => x"ffffff",
   66756 => x"ffffff",
   66757 => x"ffffff",
   66758 => x"ffffff",
   66759 => x"ffffff",
   66760 => x"ffffff",
   66761 => x"ffffff",
   66762 => x"ffffff",
   66763 => x"ffffff",
   66764 => x"ffffff",
   66765 => x"ffffff",
   66766 => x"ffffff",
   66767 => x"ffffff",
   66768 => x"ffffff",
   66769 => x"ffffff",
   66770 => x"ffffff",
   66771 => x"ffffff",
   66772 => x"ffffff",
   66773 => x"ffffff",
   66774 => x"ffffff",
   66775 => x"ffffff",
   66776 => x"ffffff",
   66777 => x"ffffff",
   66778 => x"ffffff",
   66779 => x"ffffff",
   66780 => x"ffffff",
   66781 => x"ffffff",
   66782 => x"ffffff",
   66783 => x"ffffff",
   66784 => x"ffffff",
   66785 => x"ffffff",
   66786 => x"ffffff",
   66787 => x"ffffff",
   66788 => x"ffffff",
   66789 => x"ffffff",
   66790 => x"ffffff",
   66791 => x"ffffff",
   66792 => x"ffffff",
   66793 => x"ffffff",
   66794 => x"ffffff",
   66795 => x"ffffff",
   66796 => x"ffffff",
   66797 => x"ffffff",
   66798 => x"ffffff",
   66799 => x"ffffff",
   66800 => x"ffffff",
   66801 => x"ffffff",
   66802 => x"ffffff",
   66803 => x"ffffff",
   66804 => x"ffffff",
   66805 => x"ffffff",
   66806 => x"ffffff",
   66807 => x"ffffff",
   66808 => x"ffffff",
   66809 => x"ffffff",
   66810 => x"ffffff",
   66811 => x"ffffff",
   66812 => x"ffffff",
   66813 => x"ffffff",
   66814 => x"ffffff",
   66815 => x"ffffff",
   66816 => x"ffffff",
   66817 => x"ffffff",
   66818 => x"ffffff",
   66819 => x"ffffff",
   66820 => x"ffffff",
   66821 => x"ffffff",
   66822 => x"ffffff",
   66823 => x"ffffff",
   66824 => x"ffffff",
   66825 => x"ffffff",
   66826 => x"ffffff",
   66827 => x"ffffff",
   66828 => x"ffffff",
   66829 => x"ffffff",
   66830 => x"ffffff",
   66831 => x"ffffff",
   66832 => x"ffffff",
   66833 => x"ffffff",
   66834 => x"ffffff",
   66835 => x"ffffff",
   66836 => x"ffffff",
   66837 => x"ffffff",
   66838 => x"ffffff",
   66839 => x"ffffff",
   66840 => x"ffffff",
   66841 => x"ffffff",
   66842 => x"ffffff",
   66843 => x"ffffff",
   66844 => x"ffffff",
   66845 => x"ffffff",
   66846 => x"ffffff",
   66847 => x"ffffff",
   66848 => x"ffffff",
   66849 => x"ffffff",
   66850 => x"ffffff",
   66851 => x"ffffff",
   66852 => x"ffffff",
   66853 => x"ffffff",
   66854 => x"ffffff",
   66855 => x"ffffff",
   66856 => x"ffffff",
   66857 => x"ffffff",
   66858 => x"ffffff",
   66859 => x"ffffff",
   66860 => x"ffffff",
   66861 => x"ffffff",
   66862 => x"ffffff",
   66863 => x"ffffff",
   66864 => x"ffffff",
   66865 => x"ffffff",
   66866 => x"ffffff",
   66867 => x"ffffff",
   66868 => x"ffffff",
   66869 => x"ffffff",
   66870 => x"ffffff",
   66871 => x"ffffff",
   66872 => x"ffffff",
   66873 => x"ffffff",
   66874 => x"ffffff",
   66875 => x"ffffff",
   66876 => x"ffffff",
   66877 => x"ffffff",
   66878 => x"ffffff",
   66879 => x"ffffff",
   66880 => x"ffffff",
   66881 => x"ffffff",
   66882 => x"ffffff",
   66883 => x"ffffff",
   66884 => x"ffffff",
   66885 => x"ffffff",
   66886 => x"ffffff",
   66887 => x"ffffff",
   66888 => x"ffffff",
   66889 => x"ffffff",
   66890 => x"ffffff",
   66891 => x"ffffff",
   66892 => x"ffffff",
   66893 => x"ffffff",
   66894 => x"ffffff",
   66895 => x"ffffff",
   66896 => x"ffffff",
   66897 => x"ffffff",
   66898 => x"ffffff",
   66899 => x"ffffff",
   66900 => x"ffffff",
   66901 => x"ffffff",
   66902 => x"ffffff",
   66903 => x"ffffff",
   66904 => x"ffffff",
   66905 => x"ffffff",
   66906 => x"ffffff",
   66907 => x"ffffff",
   66908 => x"ffffff",
   66909 => x"ffffff",
   66910 => x"ffffff",
   66911 => x"ffffff",
   66912 => x"ffffff",
   66913 => x"ffffff",
   66914 => x"ffffff",
   66915 => x"ffffff",
   66916 => x"ffffff",
   66917 => x"ffffff",
   66918 => x"ffffff",
   66919 => x"ffffff",
   66920 => x"ffffff",
   66921 => x"ffffff",
   66922 => x"ffffff",
   66923 => x"ffffff",
   66924 => x"ffffff",
   66925 => x"ffffff",
   66926 => x"ffffff",
   66927 => x"ffffff",
   66928 => x"ffffff",
   66929 => x"ffffff",
   66930 => x"ffffff",
   66931 => x"ffffff",
   66932 => x"ffffff",
   66933 => x"ffffff",
   66934 => x"ffffff",
   66935 => x"ffffff",
   66936 => x"ffffff",
   66937 => x"ffffff",
   66938 => x"ffffff",
   66939 => x"ffffff",
   66940 => x"ffffff",
   66941 => x"ffffff",
   66942 => x"ffffff",
   66943 => x"ffffff",
   66944 => x"ffffff",
   66945 => x"ffffff",
   66946 => x"ffffff",
   66947 => x"ffffff",
   66948 => x"ffffff",
   66949 => x"ffffff",
   66950 => x"ffffff",
   66951 => x"ffffff",
   66952 => x"ffffff",
   66953 => x"ffffff",
   66954 => x"ffffff",
   66955 => x"ffffff",
   66956 => x"ffffff",
   66957 => x"ffffff",
   66958 => x"ffffff",
   66959 => x"ffffff",
   66960 => x"ffffff",
   66961 => x"ffffff",
   66962 => x"ffffff",
   66963 => x"ffffff",
   66964 => x"ffffff",
   66965 => x"ffffff",
   66966 => x"ffffff",
   66967 => x"ffffff",
   66968 => x"ffffff",
   66969 => x"ffffff",
   66970 => x"ffffff",
   66971 => x"ffffff",
   66972 => x"ffffff",
   66973 => x"ffffff",
   66974 => x"ffffff",
   66975 => x"ffffff",
   66976 => x"ffffff",
   66977 => x"ffffff",
   66978 => x"ffffff",
   66979 => x"ffffff",
   66980 => x"ffffff",
   66981 => x"ffffff",
   66982 => x"ffffff",
   66983 => x"ffffff",
   66984 => x"ffffff",
   66985 => x"ffffff",
   66986 => x"ffffff",
   66987 => x"ffffff",
   66988 => x"ffffff",
   66989 => x"ffffff",
   66990 => x"ffffff",
   66991 => x"ffffff",
   66992 => x"ffffff",
   66993 => x"ffffff",
   66994 => x"ffffff",
   66995 => x"ffffff",
   66996 => x"ffffff",
   66997 => x"ffffff",
   66998 => x"ffffff",
   66999 => x"ffffff",
   67000 => x"ffffff",
   67001 => x"ffffff",
   67002 => x"ffffff",
   67003 => x"ffffff",
   67004 => x"ffffff",
   67005 => x"ffffff",
   67006 => x"ffffff",
   67007 => x"ffffff",
   67008 => x"ffffff",
   67009 => x"ffffff",
   67010 => x"ffffff",
   67011 => x"ffffff",
   67012 => x"ffffff",
   67013 => x"ffffff",
   67014 => x"ffffff",
   67015 => x"ffffff",
   67016 => x"ffffff",
   67017 => x"ffffff",
   67018 => x"ffffff",
   67019 => x"ffffff",
   67020 => x"ffffff",
   67021 => x"ffffff",
   67022 => x"ffffff",
   67023 => x"ffffff",
   67024 => x"ffffff",
   67025 => x"ffffff",
   67026 => x"ffffff",
   67027 => x"ffffff",
   67028 => x"ffffff",
   67029 => x"ffffff",
   67030 => x"ffffff",
   67031 => x"ffffff",
   67032 => x"ffffff",
   67033 => x"ffffff",
   67034 => x"ffffff",
   67035 => x"ffffff",
   67036 => x"ffffff",
   67037 => x"ffffff",
   67038 => x"ffffff",
   67039 => x"ffffff",
   67040 => x"ffffff",
   67041 => x"ffffff",
   67042 => x"ffffff",
   67043 => x"ffffff",
   67044 => x"ffffff",
   67045 => x"ffffff",
   67046 => x"ffffff",
   67047 => x"ffffff",
   67048 => x"ffffff",
   67049 => x"ffffff",
   67050 => x"ffffff",
   67051 => x"ffffff",
   67052 => x"ffffff",
   67053 => x"ffffff",
   67054 => x"ffffff",
   67055 => x"ffffff",
   67056 => x"ffffff",
   67057 => x"ffffff",
   67058 => x"ffffff",
   67059 => x"ffffff",
   67060 => x"ffffff",
   67061 => x"ffffff",
   67062 => x"ffffff",
   67063 => x"ffffff",
   67064 => x"ffffff",
   67065 => x"ffffff",
   67066 => x"ffffff",
   67067 => x"ffffff",
   67068 => x"ffffff",
   67069 => x"ffffff",
   67070 => x"ffffff",
   67071 => x"ffffff",
   67072 => x"ffffff",
   67073 => x"ffffff",
   67074 => x"ffffff",
   67075 => x"ffffff",
   67076 => x"ffffff",
   67077 => x"ffffff",
   67078 => x"ffffff",
   67079 => x"ffffff",
   67080 => x"ffffff",
   67081 => x"ffffff",
   67082 => x"ffffff",
   67083 => x"ffffff",
   67084 => x"ffffff",
   67085 => x"ffffff",
   67086 => x"ffffff",
   67087 => x"ffffff",
   67088 => x"ffffff",
   67089 => x"ffffff",
   67090 => x"ffffff",
   67091 => x"ffffff",
   67092 => x"ffffff",
   67093 => x"ffffff",
   67094 => x"ffffff",
   67095 => x"ffffff",
   67096 => x"ffffff",
   67097 => x"ffffff",
   67098 => x"ffffff",
   67099 => x"ffffff",
   67100 => x"ffffff",
   67101 => x"ffffff",
   67102 => x"ffffff",
   67103 => x"ffffff",
   67104 => x"ffffff",
   67105 => x"ffffff",
   67106 => x"ffffff",
   67107 => x"ffffff",
   67108 => x"ffffff",
   67109 => x"ffffff",
   67110 => x"ffffff",
   67111 => x"ffffff",
   67112 => x"ffffff",
   67113 => x"ffffff",
   67114 => x"ffffff",
   67115 => x"ffffff",
   67116 => x"ffffff",
   67117 => x"ffffff",
   67118 => x"ffffff",
   67119 => x"ffffff",
   67120 => x"ffffff",
   67121 => x"ffffff",
   67122 => x"ffffff",
   67123 => x"ffffff",
   67124 => x"ffffff",
   67125 => x"ffffff",
   67126 => x"ffffff",
   67127 => x"ffffff",
   67128 => x"ffffff",
   67129 => x"ffffff",
   67130 => x"ffffff",
   67131 => x"ffffff",
   67132 => x"ffffff",
   67133 => x"ffffff",
   67134 => x"ffffff",
   67135 => x"ffffff",
   67136 => x"ffffff",
   67137 => x"ffffff",
   67138 => x"ffffff",
   67139 => x"ffffff",
   67140 => x"ffffff",
   67141 => x"ffffff",
   67142 => x"ffffff",
   67143 => x"ffffff",
   67144 => x"ffffff",
   67145 => x"ffffff",
   67146 => x"ffffff",
   67147 => x"ffffff",
   67148 => x"ffffff",
   67149 => x"ffffff",
   67150 => x"ffffff",
   67151 => x"ffffff",
   67152 => x"ffffff",
   67153 => x"ffffff",
   67154 => x"ffffff",
   67155 => x"ffffff",
   67156 => x"ffffff",
   67157 => x"ffffff",
   67158 => x"ffffff",
   67159 => x"ffffff",
   67160 => x"ffffff",
   67161 => x"ffffff",
   67162 => x"ffffff",
   67163 => x"ffffff",
   67164 => x"ffffff",
   67165 => x"ffffff",
   67166 => x"ffffff",
   67167 => x"ffffff",
   67168 => x"ffffff",
   67169 => x"ffffff",
   67170 => x"ffffff",
   67171 => x"ffffff",
   67172 => x"ffffff",
   67173 => x"ffffff",
   67174 => x"ffffff",
   67175 => x"ffffff",
   67176 => x"ffffff",
   67177 => x"ffffff",
   67178 => x"ffffff",
   67179 => x"ffffff",
   67180 => x"ffffff",
   67181 => x"ffffff",
   67182 => x"ffffff",
   67183 => x"ffffff",
   67184 => x"ffffff",
   67185 => x"ffffff",
   67186 => x"ffffff",
   67187 => x"ffffff",
   67188 => x"ffffff",
   67189 => x"ffffff",
   67190 => x"ffffff",
   67191 => x"ffffff",
   67192 => x"ffffff",
   67193 => x"ffffff",
   67194 => x"ffffff",
   67195 => x"ffffff",
   67196 => x"ffffff",
   67197 => x"ffffff",
   67198 => x"ffffff",
   67199 => x"ffffff",
   67200 => x"ffffff",
   67201 => x"ffffff",
   67202 => x"ffffff",
   67203 => x"ffffff",
   67204 => x"ffffff",
   67205 => x"ffffff",
   67206 => x"ffffff",
   67207 => x"ffffff",
   67208 => x"ffffff",
   67209 => x"ffffff",
   67210 => x"ffffff",
   67211 => x"ffffff",
   67212 => x"ffffff",
   67213 => x"ffffff",
   67214 => x"ffffff",
   67215 => x"ffffff",
   67216 => x"ffffff",
   67217 => x"ffffff",
   67218 => x"ffffff",
   67219 => x"ffffff",
   67220 => x"ffffff",
   67221 => x"ffffff",
   67222 => x"ffffff",
   67223 => x"ffffff",
   67224 => x"ffffff",
   67225 => x"ffffff",
   67226 => x"ffffff",
   67227 => x"ffffff",
   67228 => x"ffffff",
   67229 => x"ffffff",
   67230 => x"ffffff",
   67231 => x"ffffff",
   67232 => x"ffffff",
   67233 => x"ffffff",
   67234 => x"ffffff",
   67235 => x"ffffff",
   67236 => x"ffffff",
   67237 => x"ffffff",
   67238 => x"ffffff",
   67239 => x"ffffff",
   67240 => x"ffffff",
   67241 => x"ffffff",
   67242 => x"ffffff",
   67243 => x"ffffff",
   67244 => x"ffffff",
   67245 => x"ffffff",
   67246 => x"ffffff",
   67247 => x"ffffff",
   67248 => x"ffffff",
   67249 => x"ffffff",
   67250 => x"ffffff",
   67251 => x"ffffff",
   67252 => x"ffffff",
   67253 => x"ffffff",
   67254 => x"ffffff",
   67255 => x"ffffff",
   67256 => x"ffffff",
   67257 => x"ffffff",
   67258 => x"ffffff",
   67259 => x"ffffff",
   67260 => x"ffffff",
   67261 => x"ffffff",
   67262 => x"ffffff",
   67263 => x"ffffff",
   67264 => x"ffffff",
   67265 => x"ffffff",
   67266 => x"ffffff",
   67267 => x"ffffff",
   67268 => x"ffffff",
   67269 => x"ffffff",
   67270 => x"ffffff",
   67271 => x"ffffff",
   67272 => x"ffffff",
   67273 => x"ffffff",
   67274 => x"ffffff",
   67275 => x"ffffff",
   67276 => x"ffffff",
   67277 => x"ffffff",
   67278 => x"ffffff",
   67279 => x"ffffff",
   67280 => x"ffffff",
   67281 => x"ffffff",
   67282 => x"ffffff",
   67283 => x"ffffff",
   67284 => x"ffffff",
   67285 => x"ffffff",
   67286 => x"ffffff",
   67287 => x"ffffff",
   67288 => x"ffffff",
   67289 => x"ffffff",
   67290 => x"ffffff",
   67291 => x"ffffff",
   67292 => x"ffffff",
   67293 => x"ffffff",
   67294 => x"ffffff",
   67295 => x"ffffff",
   67296 => x"ffffff",
   67297 => x"ffffff",
   67298 => x"ffffff",
   67299 => x"ffffff",
   67300 => x"ffffff",
   67301 => x"ffffff",
   67302 => x"ffffff",
   67303 => x"ffffff",
   67304 => x"ffffff",
   67305 => x"ffffff",
   67306 => x"ffffff",
   67307 => x"ffffff",
   67308 => x"ffffff",
   67309 => x"ffffff",
   67310 => x"ffffff",
   67311 => x"ffffff",
   67312 => x"ffffff",
   67313 => x"ffffff",
   67314 => x"ffffff",
   67315 => x"ffffff",
   67316 => x"ffffff",
   67317 => x"ffffff",
   67318 => x"ffffff",
   67319 => x"ffffff",
   67320 => x"ffffff",
   67321 => x"ffffff",
   67322 => x"ffffff",
   67323 => x"ffffff",
   67324 => x"ffffff",
   67325 => x"ffffff",
   67326 => x"ffffff",
   67327 => x"ffffff",
   67328 => x"ffffff",
   67329 => x"ffffff",
   67330 => x"ffffff",
   67331 => x"ffffff",
   67332 => x"ffffff",
   67333 => x"ffffff",
   67334 => x"ffffff",
   67335 => x"ffffff",
   67336 => x"ffffff",
   67337 => x"ffffff",
   67338 => x"ffffff",
   67339 => x"ffffff",
   67340 => x"ffffff",
   67341 => x"ffffff",
   67342 => x"ffffff",
   67343 => x"ffffff",
   67344 => x"ffffff",
   67345 => x"ffffff",
   67346 => x"ffffff",
   67347 => x"ffffff",
   67348 => x"ffffff",
   67349 => x"ffffff",
   67350 => x"ffffff",
   67351 => x"ffffff",
   67352 => x"ffffff",
   67353 => x"ffffff",
   67354 => x"ffffff",
   67355 => x"ffffff",
   67356 => x"ffffff",
   67357 => x"ffffff",
   67358 => x"ffffff",
   67359 => x"ffffff",
   67360 => x"ffffff",
   67361 => x"ffffff",
   67362 => x"ffffff",
   67363 => x"ffffff",
   67364 => x"ffffff",
   67365 => x"ffffff",
   67366 => x"ffffff",
   67367 => x"ffffff",
   67368 => x"ffffff",
   67369 => x"ffffff",
   67370 => x"ffffff",
   67371 => x"ffffff",
   67372 => x"ffffff",
   67373 => x"ffffff",
   67374 => x"ffffff",
   67375 => x"ffffff",
   67376 => x"ffffff",
   67377 => x"ffffff",
   67378 => x"ffffff",
   67379 => x"ffffff",
   67380 => x"ffffff",
   67381 => x"ffffff",
   67382 => x"ffffff",
   67383 => x"ffffff",
   67384 => x"ffffff",
   67385 => x"ffffff",
   67386 => x"ffffff",
   67387 => x"ffffff",
   67388 => x"ffffff",
   67389 => x"ffffff",
   67390 => x"ffffff",
   67391 => x"ffffff",
   67392 => x"ffffff",
   67393 => x"ffffff",
   67394 => x"ffffff",
   67395 => x"ffffff",
   67396 => x"ffffff",
   67397 => x"ffffff",
   67398 => x"ffffff",
   67399 => x"ffffff",
   67400 => x"ffffff",
   67401 => x"ffffff",
   67402 => x"ffffff",
   67403 => x"ffffff",
   67404 => x"ffffff",
   67405 => x"ffffff",
   67406 => x"ffffff",
   67407 => x"ffffff",
   67408 => x"ffffff",
   67409 => x"ffffff",
   67410 => x"ffffff",
   67411 => x"ffffff",
   67412 => x"ffffff",
   67413 => x"ffffff",
   67414 => x"ffffff",
   67415 => x"ffffff",
   67416 => x"ffffff",
   67417 => x"ffffff",
   67418 => x"ffffff",
   67419 => x"ffffff",
   67420 => x"ffffff",
   67421 => x"ffffff",
   67422 => x"ffffff",
   67423 => x"ffffff",
   67424 => x"ffffff",
   67425 => x"ffffff",
   67426 => x"ffffff",
   67427 => x"ffffff",
   67428 => x"ffffff",
   67429 => x"ffffff",
   67430 => x"ffffff",
   67431 => x"ffffff",
   67432 => x"ffffff",
   67433 => x"ffffff",
   67434 => x"ffffff",
   67435 => x"ffffff",
   67436 => x"ffffff",
   67437 => x"ffffff",
   67438 => x"ffffff",
   67439 => x"ffffff",
   67440 => x"ffffff",
   67441 => x"ffffff",
   67442 => x"ffffff",
   67443 => x"ffffff",
   67444 => x"ffffff",
   67445 => x"ffffff",
   67446 => x"ffffff",
   67447 => x"ffffff",
   67448 => x"ffffff",
   67449 => x"ffffff",
   67450 => x"ffffff",
   67451 => x"ffffff",
   67452 => x"ffffff",
   67453 => x"ffffff",
   67454 => x"ffffff",
   67455 => x"ffffff",
   67456 => x"ffffff",
   67457 => x"ffffff",
   67458 => x"ffffff",
   67459 => x"ffffff",
   67460 => x"ffffff",
   67461 => x"ffffff",
   67462 => x"ffffff",
   67463 => x"ffffff",
   67464 => x"ffffff",
   67465 => x"ffffff",
   67466 => x"ffffff",
   67467 => x"ffffff",
   67468 => x"ffffff",
   67469 => x"ffffff",
   67470 => x"ffffff",
   67471 => x"ffffff",
   67472 => x"ffffff",
   67473 => x"ffffff",
   67474 => x"ffffff",
   67475 => x"ffffff",
   67476 => x"ffffff",
   67477 => x"ffffff",
   67478 => x"ffffff",
   67479 => x"ffffff",
   67480 => x"ffffff",
   67481 => x"ffffff",
   67482 => x"ffffff",
   67483 => x"ffffff",
   67484 => x"ffffff",
   67485 => x"ffffff",
   67486 => x"ffffff",
   67487 => x"ffffff",
   67488 => x"ffffff",
   67489 => x"ffffff",
   67490 => x"ffffff",
   67491 => x"ffffff",
   67492 => x"ffffff",
   67493 => x"ffffff",
   67494 => x"ffffff",
   67495 => x"ffffff",
   67496 => x"ffffff",
   67497 => x"ffffff",
   67498 => x"ffffff",
   67499 => x"ffffff",
   67500 => x"ffffff",
   67501 => x"ffffff",
   67502 => x"ffffff",
   67503 => x"ffffff",
   67504 => x"ffffff",
   67505 => x"ffffff",
   67506 => x"ffffff",
   67507 => x"ffffff",
   67508 => x"ffffff",
   67509 => x"ffffff",
   67510 => x"ffffff",
   67511 => x"ffffff",
   67512 => x"ffffff",
   67513 => x"ffffff",
   67514 => x"ffffff",
   67515 => x"ffffff",
   67516 => x"ffffff",
   67517 => x"ffffff",
   67518 => x"ffffff",
   67519 => x"ffffff",
   67520 => x"ffffff",
   67521 => x"ffffff",
   67522 => x"ffffff",
   67523 => x"ffffff",
   67524 => x"ffffff",
   67525 => x"ffffff",
   67526 => x"ffffff",
   67527 => x"ffffff",
   67528 => x"ffffff",
   67529 => x"ffffff",
   67530 => x"ffffff",
   67531 => x"ffffff",
   67532 => x"ffffff",
   67533 => x"ffffff",
   67534 => x"ffffff",
   67535 => x"ffffff",
   67536 => x"ffffff",
   67537 => x"ffffff",
   67538 => x"ffffff",
   67539 => x"ffffff",
   67540 => x"ffffff",
   67541 => x"ffffff",
   67542 => x"ffffff",
   67543 => x"ffffff",
   67544 => x"ffffff",
   67545 => x"ffffff",
   67546 => x"ffffff",
   67547 => x"ffffff",
   67548 => x"ffffff",
   67549 => x"ffffff",
   67550 => x"ffffff",
   67551 => x"ffffff",
   67552 => x"ffffff",
   67553 => x"ffffff",
   67554 => x"ffffff",
   67555 => x"ffffff",
   67556 => x"ffffff",
   67557 => x"ffffff",
   67558 => x"ffffff",
   67559 => x"ffffff",
   67560 => x"ffffff",
   67561 => x"ffffff",
   67562 => x"ffffff",
   67563 => x"ffffff",
   67564 => x"ffffff",
   67565 => x"ffffff",
   67566 => x"ffffff",
   67567 => x"ffffff",
   67568 => x"ffffff",
   67569 => x"ffffff",
   67570 => x"ffffff",
   67571 => x"ffffff",
   67572 => x"ffffff",
   67573 => x"ffffff",
   67574 => x"ffffff",
   67575 => x"ffffff",
   67576 => x"ffffff",
   67577 => x"ffffff",
   67578 => x"ffffff",
   67579 => x"ffffff",
   67580 => x"ffffff",
   67581 => x"ffffff",
   67582 => x"ffffff",
   67583 => x"ffffff",
   67584 => x"ffffff",
   67585 => x"ffffff",
   67586 => x"ffffff",
   67587 => x"ffffff",
   67588 => x"ffffff",
   67589 => x"ffffff",
   67590 => x"ffffff",
   67591 => x"ffffff",
   67592 => x"ffffff",
   67593 => x"ffffff",
   67594 => x"ffffff",
   67595 => x"ffffff",
   67596 => x"ffffff",
   67597 => x"ffffff",
   67598 => x"ffffff",
   67599 => x"ffffff",
   67600 => x"ffffff",
   67601 => x"ffffff",
   67602 => x"ffffff",
   67603 => x"ffffff",
   67604 => x"ffffff",
   67605 => x"ffffff",
   67606 => x"ffffff",
   67607 => x"ffffff",
   67608 => x"ffffff",
   67609 => x"ffffff",
   67610 => x"ffffff",
   67611 => x"ffffff",
   67612 => x"ffffff",
   67613 => x"ffffff",
   67614 => x"ffffff",
   67615 => x"ffffff",
   67616 => x"ffffff",
   67617 => x"ffffff",
   67618 => x"ffffff",
   67619 => x"ffffff",
   67620 => x"ffffff",
   67621 => x"ffffff",
   67622 => x"ffffff",
   67623 => x"ffffff",
   67624 => x"ffffff",
   67625 => x"ffffff",
   67626 => x"ffffff",
   67627 => x"ffffff",
   67628 => x"ffffff",
   67629 => x"ffffff",
   67630 => x"ffffff",
   67631 => x"ffffff",
   67632 => x"ffffff",
   67633 => x"ffffff",
   67634 => x"ffffff",
   67635 => x"ffffff",
   67636 => x"ffffff",
   67637 => x"ffffff",
   67638 => x"ffffff",
   67639 => x"ffffff",
   67640 => x"ffffff",
   67641 => x"ffffff",
   67642 => x"ffffff",
   67643 => x"ffffff",
   67644 => x"ffffff",
   67645 => x"ffffff",
   67646 => x"ffffff",
   67647 => x"ffffff",
   67648 => x"ffffff",
   67649 => x"ffffff",
   67650 => x"ffffff",
   67651 => x"ffffff",
   67652 => x"ffffff",
   67653 => x"ffffff",
   67654 => x"ffffff",
   67655 => x"ffffff",
   67656 => x"ffffff",
   67657 => x"ffffff",
   67658 => x"ffffff",
   67659 => x"ffffff",
   67660 => x"ffffff",
   67661 => x"ffffff",
   67662 => x"ffffff",
   67663 => x"ffffff",
   67664 => x"ffffff",
   67665 => x"ffffff",
   67666 => x"ffffff",
   67667 => x"ffffff",
   67668 => x"ffffff",
   67669 => x"ffffff",
   67670 => x"ffffff",
   67671 => x"ffffff",
   67672 => x"ffffff",
   67673 => x"ffffff",
   67674 => x"ffffff",
   67675 => x"ffffff",
   67676 => x"ffffff",
   67677 => x"ffffff",
   67678 => x"ffffff",
   67679 => x"ffffff",
   67680 => x"ffffff",
   67681 => x"ffffff",
   67682 => x"ffffff",
   67683 => x"ffffff",
   67684 => x"ffffff",
   67685 => x"ffffff",
   67686 => x"ffffff",
   67687 => x"ffffff",
   67688 => x"ffffff",
   67689 => x"ffffff",
   67690 => x"ffffff",
   67691 => x"ffffff",
   67692 => x"ffffff",
   67693 => x"ffffff",
   67694 => x"ffffff",
   67695 => x"ffffff",
   67696 => x"ffffff",
   67697 => x"ffffff",
   67698 => x"ffffff",
   67699 => x"ffffff",
   67700 => x"ffffff",
   67701 => x"ffffff",
   67702 => x"ffffff",
   67703 => x"ffffff",
   67704 => x"ffffff",
   67705 => x"ffffff",
   67706 => x"ffffff",
   67707 => x"ffffff",
   67708 => x"ffffff",
   67709 => x"ffffff",
   67710 => x"ffffff",
   67711 => x"ffffff",
   67712 => x"ffffff",
   67713 => x"ffffff",
   67714 => x"ffffff",
   67715 => x"ffffff",
   67716 => x"ffffff",
   67717 => x"ffffff",
   67718 => x"ffffff",
   67719 => x"ffffff",
   67720 => x"ffffff",
   67721 => x"ffffff",
   67722 => x"ffffff",
   67723 => x"ffffff",
   67724 => x"ffffff",
   67725 => x"ffffff",
   67726 => x"ffffff",
   67727 => x"ffffff",
   67728 => x"ffffff",
   67729 => x"ffffff",
   67730 => x"ffffff",
   67731 => x"ffffff",
   67732 => x"ffffff",
   67733 => x"ffffff",
   67734 => x"ffffff",
   67735 => x"ffffff",
   67736 => x"ffffff",
   67737 => x"ffffff",
   67738 => x"ffffff",
   67739 => x"ffffff",
   67740 => x"ffffff",
   67741 => x"ffffff",
   67742 => x"ffffff",
   67743 => x"ffffff",
   67744 => x"ffffff",
   67745 => x"ffffff",
   67746 => x"ffffff",
   67747 => x"ffffff",
   67748 => x"ffffff",
   67749 => x"ffffff",
   67750 => x"ffffff",
   67751 => x"ffffff",
   67752 => x"ffffff",
   67753 => x"ffffff",
   67754 => x"ffffff",
   67755 => x"ffffff",
   67756 => x"ffffff",
   67757 => x"ffffff",
   67758 => x"ffffff",
   67759 => x"ffffff",
   67760 => x"ffffff",
   67761 => x"ffffff",
   67762 => x"ffffff",
   67763 => x"ffffff",
   67764 => x"ffffff",
   67765 => x"ffffff",
   67766 => x"ffffff",
   67767 => x"ffffff",
   67768 => x"ffffff",
   67769 => x"ffffff",
   67770 => x"ffffff",
   67771 => x"ffffff",
   67772 => x"ffffff",
   67773 => x"ffffff",
   67774 => x"ffffff",
   67775 => x"ffffff",
   67776 => x"ffffff",
   67777 => x"ffffff",
   67778 => x"ffffff",
   67779 => x"ffffff",
   67780 => x"ffffff",
   67781 => x"ffffff",
   67782 => x"ffffff",
   67783 => x"ffffff",
   67784 => x"ffffff",
   67785 => x"ffffff",
   67786 => x"ffffff",
   67787 => x"ffffff",
   67788 => x"ffffff",
   67789 => x"ffffff",
   67790 => x"ffffff",
   67791 => x"ffffff",
   67792 => x"ffffff",
   67793 => x"ffffff",
   67794 => x"ffffff",
   67795 => x"ffffff",
   67796 => x"ffffff",
   67797 => x"ffffff",
   67798 => x"ffffff",
   67799 => x"ffffff",
   67800 => x"ffffff",
   67801 => x"ffffff",
   67802 => x"ffffff",
   67803 => x"ffffff",
   67804 => x"ffffff",
   67805 => x"ffffff",
   67806 => x"ffffff",
   67807 => x"ffffff",
   67808 => x"ffffff",
   67809 => x"ffffff",
   67810 => x"ffffff",
   67811 => x"ffffff",
   67812 => x"ffffff",
   67813 => x"ffffff",
   67814 => x"ffffff",
   67815 => x"ffffff",
   67816 => x"ffffff",
   67817 => x"ffffff",
   67818 => x"ffffff",
   67819 => x"ffffff",
   67820 => x"ffffff",
   67821 => x"ffffff",
   67822 => x"ffffff",
   67823 => x"ffffff",
   67824 => x"ffffff",
   67825 => x"ffffff",
   67826 => x"ffffff",
   67827 => x"ffffff",
   67828 => x"ffffff",
   67829 => x"ffffff",
   67830 => x"ffffff",
   67831 => x"ffffff",
   67832 => x"ffffff",
   67833 => x"ffffff",
   67834 => x"ffffff",
   67835 => x"ffffff",
   67836 => x"ffffff",
   67837 => x"ffffff",
   67838 => x"ffffff",
   67839 => x"ffffff",
   67840 => x"ffffff",
   67841 => x"ffffff",
   67842 => x"ffffff",
   67843 => x"ffffff",
   67844 => x"ffffff",
   67845 => x"ffffff",
   67846 => x"ffffff",
   67847 => x"ffffff",
   67848 => x"ffffff",
   67849 => x"ffffff",
   67850 => x"ffffff",
   67851 => x"ffffff",
   67852 => x"ffffff",
   67853 => x"ffffff",
   67854 => x"ffffff",
   67855 => x"ffffff",
   67856 => x"ffffff",
   67857 => x"ffffff",
   67858 => x"ffffff",
   67859 => x"ffffff",
   67860 => x"ffffff",
   67861 => x"ffffff",
   67862 => x"ffffff",
   67863 => x"ffffff",
   67864 => x"ffffff",
   67865 => x"ffffff",
   67866 => x"ffffff",
   67867 => x"ffffff",
   67868 => x"ffffff",
   67869 => x"ffffff",
   67870 => x"ffffff",
   67871 => x"ffffff",
   67872 => x"ffffff",
   67873 => x"ffffff",
   67874 => x"ffffff",
   67875 => x"ffffff",
   67876 => x"ffffff",
   67877 => x"ffffff",
   67878 => x"ffffff",
   67879 => x"ffffff",
   67880 => x"ffffff",
   67881 => x"ffffff",
   67882 => x"ffffff",
   67883 => x"ffffff",
   67884 => x"ffffff",
   67885 => x"ffffff",
   67886 => x"ffffff",
   67887 => x"ffffff",
   67888 => x"ffffff",
   67889 => x"ffffff",
   67890 => x"ffffff",
   67891 => x"ffffff",
   67892 => x"ffffff",
   67893 => x"ffffff",
   67894 => x"ffffff",
   67895 => x"ffffff",
   67896 => x"ffffff",
   67897 => x"ffffff",
   67898 => x"ffffff",
   67899 => x"ffffff",
   67900 => x"ffffff",
   67901 => x"ffffff",
   67902 => x"ffffff",
   67903 => x"ffffff",
   67904 => x"ffffff",
   67905 => x"ffffff",
   67906 => x"ffffff",
   67907 => x"ffffff",
   67908 => x"ffffff",
   67909 => x"ffffff",
   67910 => x"ffffff",
   67911 => x"ffffff",
   67912 => x"ffffff",
   67913 => x"ffffff",
   67914 => x"ffffff",
   67915 => x"ffffff",
   67916 => x"ffffff",
   67917 => x"ffffff",
   67918 => x"ffffff",
   67919 => x"ffffff",
   67920 => x"ffffff",
   67921 => x"ffffff",
   67922 => x"ffffff",
   67923 => x"ffffff",
   67924 => x"ffffff",
   67925 => x"ffffff",
   67926 => x"ffffff",
   67927 => x"ffffff",
   67928 => x"ffffff",
   67929 => x"ffffff",
   67930 => x"ffffff",
   67931 => x"ffffff",
   67932 => x"ffffff",
   67933 => x"ffffff",
   67934 => x"ffffff",
   67935 => x"ffffff",
   67936 => x"ffffff",
   67937 => x"ffffff",
   67938 => x"ffffff",
   67939 => x"ffffff",
   67940 => x"ffffff",
   67941 => x"ffffff",
   67942 => x"ffffff",
   67943 => x"ffffff",
   67944 => x"ffffff",
   67945 => x"ffffff",
   67946 => x"ffffff",
   67947 => x"ffffff",
   67948 => x"ffffff",
   67949 => x"ffffff",
   67950 => x"ffffff",
   67951 => x"ffffff",
   67952 => x"ffffff",
   67953 => x"ffffff",
   67954 => x"ffffff",
   67955 => x"ffffff",
   67956 => x"ffffff",
   67957 => x"ffffff",
   67958 => x"ffffff",
   67959 => x"ffffff",
   67960 => x"ffffff",
   67961 => x"ffffff",
   67962 => x"ffffff",
   67963 => x"ffffff",
   67964 => x"ffffff",
   67965 => x"ffffff",
   67966 => x"ffffff",
   67967 => x"ffffff",
   67968 => x"ffffff",
   67969 => x"ffffff",
   67970 => x"ffffff",
   67971 => x"ffffff",
   67972 => x"ffffff",
   67973 => x"ffffff",
   67974 => x"ffffff",
   67975 => x"ffffff",
   67976 => x"ffffff",
   67977 => x"ffffff",
   67978 => x"ffffff",
   67979 => x"ffffff",
   67980 => x"ffffff",
   67981 => x"ffffff",
   67982 => x"ffffff",
   67983 => x"ffffff",
   67984 => x"ffffff",
   67985 => x"ffffff",
   67986 => x"ffffff",
   67987 => x"ffffff",
   67988 => x"ffffff",
   67989 => x"ffffff",
   67990 => x"ffffff",
   67991 => x"ffffff",
   67992 => x"ffffff",
   67993 => x"ffffff",
   67994 => x"ffffff",
   67995 => x"ffffff",
   67996 => x"ffffff",
   67997 => x"ffffff",
   67998 => x"ffffff",
   67999 => x"ffffff",
   68000 => x"ffffff",
   68001 => x"ffffff",
   68002 => x"ffffff",
   68003 => x"ffffff",
   68004 => x"ffffff",
   68005 => x"ffffff",
   68006 => x"ffffff",
   68007 => x"ffffff",
   68008 => x"ffffff",
   68009 => x"ffffff",
   68010 => x"ffffff",
   68011 => x"ffffff",
   68012 => x"ffffff",
   68013 => x"ffffff",
   68014 => x"ffffff",
   68015 => x"ffffff",
   68016 => x"ffffff",
   68017 => x"ffffff",
   68018 => x"ffffff",
   68019 => x"ffffff",
   68020 => x"ffffff",
   68021 => x"ffffff",
   68022 => x"ffffff",
   68023 => x"ffffff",
   68024 => x"ffffff",
   68025 => x"ffffff",
   68026 => x"ffffff",
   68027 => x"ffffff",
   68028 => x"ffffff",
   68029 => x"ffffff",
   68030 => x"ffffff",
   68031 => x"ffffff",
   68032 => x"ffffff",
   68033 => x"ffffff",
   68034 => x"ffffff",
   68035 => x"ffffff",
   68036 => x"ffffff",
   68037 => x"ffffff",
   68038 => x"ffffff",
   68039 => x"ffffff",
   68040 => x"ffffff",
   68041 => x"ffffff",
   68042 => x"ffffff",
   68043 => x"ffffff",
   68044 => x"ffffff",
   68045 => x"ffffff",
   68046 => x"ffffff",
   68047 => x"ffffff",
   68048 => x"ffffff",
   68049 => x"ffffff",
   68050 => x"ffffff",
   68051 => x"ffffff",
   68052 => x"ffffff",
   68053 => x"ffffff",
   68054 => x"ffffff",
   68055 => x"ffffff",
   68056 => x"ffffff",
   68057 => x"ffffff",
   68058 => x"ffffff",
   68059 => x"ffffff",
   68060 => x"ffffff",
   68061 => x"ffffff",
   68062 => x"ffffff",
   68063 => x"ffffff",
   68064 => x"ffffff",
   68065 => x"ffffff",
   68066 => x"ffffff",
   68067 => x"ffffff",
   68068 => x"ffffff",
   68069 => x"ffffff",
   68070 => x"ffffff",
   68071 => x"ffffff",
   68072 => x"ffffff",
   68073 => x"ffffff",
   68074 => x"ffffff",
   68075 => x"ffffff",
   68076 => x"ffffff",
   68077 => x"ffffff",
   68078 => x"ffffff",
   68079 => x"ffffff",
   68080 => x"ffffff",
   68081 => x"ffffff",
   68082 => x"ffffff",
   68083 => x"ffffff",
   68084 => x"ffffff",
   68085 => x"ffffff",
   68086 => x"ffffff",
   68087 => x"ffffff",
   68088 => x"ffffff",
   68089 => x"ffffff",
   68090 => x"ffffff",
   68091 => x"ffffff",
   68092 => x"ffffff",
   68093 => x"ffffff",
   68094 => x"ffffff",
   68095 => x"ffffff",
   68096 => x"ffffff",
   68097 => x"ffffff",
   68098 => x"ffffff",
   68099 => x"ffffff",
   68100 => x"ffffff",
   68101 => x"ffffff",
   68102 => x"ffffff",
   68103 => x"ffffff",
   68104 => x"ffffff",
   68105 => x"ffffff",
   68106 => x"ffffff",
   68107 => x"ffffff",
   68108 => x"ffffff",
   68109 => x"ffffff",
   68110 => x"ffffff",
   68111 => x"ffffff",
   68112 => x"ffffff",
   68113 => x"ffffff",
   68114 => x"ffffff",
   68115 => x"ffffff",
   68116 => x"ffffff",
   68117 => x"ffffff",
   68118 => x"ffffff",
   68119 => x"ffffff",
   68120 => x"ffffff",
   68121 => x"ffffff",
   68122 => x"ffffff",
   68123 => x"ffffff",
   68124 => x"ffffff",
   68125 => x"ffffff",
   68126 => x"ffffff",
   68127 => x"ffffff",
   68128 => x"ffffff",
   68129 => x"ffffff",
   68130 => x"ffffff",
   68131 => x"ffffff",
   68132 => x"ffffff",
   68133 => x"ffffff",
   68134 => x"ffffff",
   68135 => x"ffffff",
   68136 => x"ffffff",
   68137 => x"ffffff",
   68138 => x"ffffff",
   68139 => x"ffffff",
   68140 => x"ffffff",
   68141 => x"ffffff",
   68142 => x"ffffff",
   68143 => x"ffffff",
   68144 => x"ffffff",
   68145 => x"ffffff",
   68146 => x"ffffff",
   68147 => x"ffffff",
   68148 => x"ffffff",
   68149 => x"ffffff",
   68150 => x"ffffff",
   68151 => x"ffffff",
   68152 => x"ffffff",
   68153 => x"ffffff",
   68154 => x"ffffff",
   68155 => x"ffffff",
   68156 => x"ffffff",
   68157 => x"ffffff",
   68158 => x"ffffff",
   68159 => x"ffffff",
   68160 => x"ffffff",
   68161 => x"ffffff",
   68162 => x"ffffff",
   68163 => x"ffffff",
   68164 => x"ffffff",
   68165 => x"ffffff",
   68166 => x"ffffff",
   68167 => x"ffffff",
   68168 => x"ffffff",
   68169 => x"ffffff",
   68170 => x"ffffff",
   68171 => x"ffffff",
   68172 => x"ffffff",
   68173 => x"ffffff",
   68174 => x"ffffff",
   68175 => x"ffffff",
   68176 => x"ffffff",
   68177 => x"ffffff",
   68178 => x"ffffff",
   68179 => x"ffffff",
   68180 => x"ffffff",
   68181 => x"ffffff",
   68182 => x"ffffff",
   68183 => x"ffffff",
   68184 => x"ffffff",
   68185 => x"ffffff",
   68186 => x"ffffff",
   68187 => x"ffffff",
   68188 => x"ffffff",
   68189 => x"ffffff",
   68190 => x"ffffff",
   68191 => x"ffffff",
   68192 => x"ffffff",
   68193 => x"ffffff",
   68194 => x"ffffff",
   68195 => x"ffffff",
   68196 => x"ffffff",
   68197 => x"ffffff",
   68198 => x"ffffff",
   68199 => x"ffffff",
   68200 => x"ffffff",
   68201 => x"ffffff",
   68202 => x"ffffff",
   68203 => x"ffffff",
   68204 => x"ffffff",
   68205 => x"ffffff",
   68206 => x"ffffff",
   68207 => x"ffffff",
   68208 => x"ffffff",
   68209 => x"ffffff",
   68210 => x"ffffff",
   68211 => x"ffffff",
   68212 => x"ffffff",
   68213 => x"ffffff",
   68214 => x"ffffff",
   68215 => x"ffffff",
   68216 => x"ffffff",
   68217 => x"ffffff",
   68218 => x"ffffff",
   68219 => x"ffffff",
   68220 => x"ffffff",
   68221 => x"ffffff",
   68222 => x"ffffff",
   68223 => x"ffffff",
   68224 => x"ffffff",
   68225 => x"ffffff",
   68226 => x"ffffff",
   68227 => x"ffffff",
   68228 => x"ffffff",
   68229 => x"ffffff",
   68230 => x"ffffff",
   68231 => x"ffffff",
   68232 => x"ffffff",
   68233 => x"ffffff",
   68234 => x"ffffff",
   68235 => x"ffffff",
   68236 => x"ffffff",
   68237 => x"ffffff",
   68238 => x"ffffff",
   68239 => x"ffffff",
   68240 => x"ffffff",
   68241 => x"ffffff",
   68242 => x"ffffff",
   68243 => x"ffffff",
   68244 => x"ffffff",
   68245 => x"ffffff",
   68246 => x"ffffff",
   68247 => x"ffffff",
   68248 => x"ffffff",
   68249 => x"ffffff",
   68250 => x"ffffff",
   68251 => x"ffffff",
   68252 => x"ffffff",
   68253 => x"ffffff",
   68254 => x"ffffff",
   68255 => x"ffffff",
   68256 => x"ffffff",
   68257 => x"ffffff",
   68258 => x"ffffff",
   68259 => x"ffffff",
   68260 => x"ffffff",
   68261 => x"ffffff",
   68262 => x"ffffff",
   68263 => x"ffffff",
   68264 => x"ffffff",
   68265 => x"ffffff",
   68266 => x"ffffff",
   68267 => x"ffffff",
   68268 => x"ffffff",
   68269 => x"ffffff",
   68270 => x"ffffff",
   68271 => x"ffffff",
   68272 => x"ffffff",
   68273 => x"ffffff",
   68274 => x"ffffff",
   68275 => x"ffffff",
   68276 => x"ffffff",
   68277 => x"ffffff",
   68278 => x"ffffff",
   68279 => x"ffffff",
   68280 => x"ffffff",
   68281 => x"ffffff",
   68282 => x"ffffff",
   68283 => x"ffffff",
   68284 => x"ffffff",
   68285 => x"ffffff",
   68286 => x"ffffff",
   68287 => x"ffffff",
   68288 => x"ffffff",
   68289 => x"ffffff",
   68290 => x"ffffff",
   68291 => x"ffffff",
   68292 => x"ffffff",
   68293 => x"ffffff",
   68294 => x"ffffff",
   68295 => x"ffffff",
   68296 => x"ffffff",
   68297 => x"ffffff",
   68298 => x"ffffff",
   68299 => x"ffffff",
   68300 => x"ffffff",
   68301 => x"ffffff",
   68302 => x"ffffff",
   68303 => x"ffffff",
   68304 => x"ffffff",
   68305 => x"ffffff",
   68306 => x"ffffff",
   68307 => x"ffffff",
   68308 => x"ffffff",
   68309 => x"ffffff",
   68310 => x"ffffff",
   68311 => x"ffffff",
   68312 => x"ffffff",
   68313 => x"ffffff",
   68314 => x"ffffff",
   68315 => x"ffffff",
   68316 => x"ffffff",
   68317 => x"ffffff",
   68318 => x"ffffff",
   68319 => x"ffffff",
   68320 => x"ffffff",
   68321 => x"ffffff",
   68322 => x"ffffff",
   68323 => x"ffffff",
   68324 => x"ffffff",
   68325 => x"ffffff",
   68326 => x"ffffff",
   68327 => x"ffffff",
   68328 => x"ffffff",
   68329 => x"ffffff",
   68330 => x"ffffff",
   68331 => x"ffffff",
   68332 => x"ffffff",
   68333 => x"ffffff",
   68334 => x"ffffff",
   68335 => x"ffffff",
   68336 => x"ffffff",
   68337 => x"ffffff",
   68338 => x"ffffff",
   68339 => x"ffffff",
   68340 => x"ffffff",
   68341 => x"ffffff",
   68342 => x"ffffff",
   68343 => x"ffffff",
   68344 => x"ffffff",
   68345 => x"ffffff",
   68346 => x"ffffff",
   68347 => x"ffffff",
   68348 => x"ffffff",
   68349 => x"ffffff",
   68350 => x"ffffff",
   68351 => x"ffffff",
   68352 => x"ffffff",
   68353 => x"ffffff",
   68354 => x"ffffff",
   68355 => x"ffffff",
   68356 => x"ffffff",
   68357 => x"ffffff",
   68358 => x"ffffff",
   68359 => x"ffffff",
   68360 => x"ffffff",
   68361 => x"ffffff",
   68362 => x"ffffff",
   68363 => x"ffffff",
   68364 => x"ffffff",
   68365 => x"ffffff",
   68366 => x"ffffff",
   68367 => x"ffffff",
   68368 => x"ffffff",
   68369 => x"ffffff",
   68370 => x"ffffff",
   68371 => x"ffffff",
   68372 => x"ffffff",
   68373 => x"ffffff",
   68374 => x"ffffff",
   68375 => x"ffffff",
   68376 => x"ffffff",
   68377 => x"ffffff",
   68378 => x"ffffff",
   68379 => x"ffffff",
   68380 => x"ffffff",
   68381 => x"ffffff",
   68382 => x"ffffff",
   68383 => x"ffffff",
   68384 => x"ffffff",
   68385 => x"ffffff",
   68386 => x"ffffff",
   68387 => x"ffffff",
   68388 => x"ffffff",
   68389 => x"ffffff",
   68390 => x"ffffff",
   68391 => x"ffffff",
   68392 => x"ffffff",
   68393 => x"ffffff",
   68394 => x"ffffff",
   68395 => x"ffffff",
   68396 => x"ffffff",
   68397 => x"ffffff",
   68398 => x"ffffff",
   68399 => x"ffffff",
   68400 => x"ffffff",
   68401 => x"ffffff",
   68402 => x"ffffff",
   68403 => x"ffffff",
   68404 => x"ffffff",
   68405 => x"ffffff",
   68406 => x"ffffff",
   68407 => x"ffffff",
   68408 => x"ffffff",
   68409 => x"ffffff",
   68410 => x"ffffff",
   68411 => x"ffffff",
   68412 => x"ffffff",
   68413 => x"ffffff",
   68414 => x"ffffff",
   68415 => x"ffffff",
   68416 => x"ffffff",
   68417 => x"ffffff",
   68418 => x"ffffff",
   68419 => x"ffffff",
   68420 => x"ffffff",
   68421 => x"ffffff",
   68422 => x"ffffff",
   68423 => x"ffffff",
   68424 => x"ffffff",
   68425 => x"ffffff",
   68426 => x"ffffff",
   68427 => x"ffffff",
   68428 => x"ffffff",
   68429 => x"ffffff",
   68430 => x"ffffff",
   68431 => x"ffffff",
   68432 => x"ffffff",
   68433 => x"ffffff",
   68434 => x"ffffff",
   68435 => x"ffffff",
   68436 => x"ffffff",
   68437 => x"ffffff",
   68438 => x"ffffff",
   68439 => x"ffffff",
   68440 => x"ffffff",
   68441 => x"ffffff",
   68442 => x"ffffff",
   68443 => x"ffffff",
   68444 => x"ffffff",
   68445 => x"ffffff",
   68446 => x"ffffff",
   68447 => x"ffffff",
   68448 => x"ffffff",
   68449 => x"ffffff",
   68450 => x"ffffff",
   68451 => x"ffffff",
   68452 => x"ffffff",
   68453 => x"ffffff",
   68454 => x"ffffff",
   68455 => x"ffffff",
   68456 => x"ffffff",
   68457 => x"ffffff",
   68458 => x"ffffff",
   68459 => x"ffffff",
   68460 => x"ffffff",
   68461 => x"ffffff",
   68462 => x"ffffff",
   68463 => x"ffffff",
   68464 => x"ffffff",
   68465 => x"ffffff",
   68466 => x"ffffff",
   68467 => x"ffffff",
   68468 => x"ffffff",
   68469 => x"ffffff",
   68470 => x"ffffff",
   68471 => x"ffffff",
   68472 => x"ffffff",
   68473 => x"ffffff",
   68474 => x"ffffff",
   68475 => x"ffffff",
   68476 => x"ffffff",
   68477 => x"ffffff",
   68478 => x"ffffff",
   68479 => x"ffffff",
   68480 => x"ffffff",
   68481 => x"ffffff",
   68482 => x"ffffff",
   68483 => x"ffffff",
   68484 => x"ffffff",
   68485 => x"ffffff",
   68486 => x"ffffff",
   68487 => x"ffffff",
   68488 => x"ffffff",
   68489 => x"ffffff",
   68490 => x"ffffff",
   68491 => x"ffffff",
   68492 => x"ffffff",
   68493 => x"ffffff",
   68494 => x"ffffff",
   68495 => x"ffffff",
   68496 => x"ffffff",
   68497 => x"ffffff",
   68498 => x"ffffff",
   68499 => x"ffffff",
   68500 => x"ffffff",
   68501 => x"ffffff",
   68502 => x"ffffff",
   68503 => x"ffffff",
   68504 => x"ffffff",
   68505 => x"ffffff",
   68506 => x"ffffff",
   68507 => x"ffffff",
   68508 => x"ffffff",
   68509 => x"ffffff",
   68510 => x"ffffff",
   68511 => x"ffffff",
   68512 => x"ffffff",
   68513 => x"ffffff",
   68514 => x"ffffff",
   68515 => x"ffffff",
   68516 => x"ffffff",
   68517 => x"ffffff",
   68518 => x"ffffff",
   68519 => x"ffffff",
   68520 => x"ffffff",
   68521 => x"ffffff",
   68522 => x"ffffff",
   68523 => x"ffffff",
   68524 => x"ffffff",
   68525 => x"ffffff",
   68526 => x"ffffff",
   68527 => x"ffffff",
   68528 => x"ffffff",
   68529 => x"ffffff",
   68530 => x"ffffff",
   68531 => x"ffffff",
   68532 => x"ffffff",
   68533 => x"ffffff",
   68534 => x"ffffff",
   68535 => x"ffffff",
   68536 => x"ffffff",
   68537 => x"ffffff",
   68538 => x"ffffff",
   68539 => x"ffffff",
   68540 => x"ffffff",
   68541 => x"ffffff",
   68542 => x"ffffff",
   68543 => x"ffffff",
   68544 => x"ffffff",
   68545 => x"ffffff",
   68546 => x"ffffff",
   68547 => x"ffffff",
   68548 => x"ffffff",
   68549 => x"ffffff",
   68550 => x"ffffff",
   68551 => x"ffffff",
   68552 => x"ffffff",
   68553 => x"ffffff",
   68554 => x"ffffff",
   68555 => x"ffffff",
   68556 => x"ffffff",
   68557 => x"ffffff",
   68558 => x"ffffff",
   68559 => x"ffffff",
   68560 => x"ffffff",
   68561 => x"ffffff",
   68562 => x"ffffff",
   68563 => x"ffffff",
   68564 => x"ffffff",
   68565 => x"ffffff",
   68566 => x"ffffff",
   68567 => x"ffffff",
   68568 => x"ffffff",
   68569 => x"ffffff",
   68570 => x"ffffff",
   68571 => x"ffffff",
   68572 => x"ffffff",
   68573 => x"ffffff",
   68574 => x"ffffff",
   68575 => x"ffffff",
   68576 => x"ffffff",
   68577 => x"ffffff",
   68578 => x"ffffff",
   68579 => x"ffffff",
   68580 => x"ffffff",
   68581 => x"ffffff",
   68582 => x"ffffff",
   68583 => x"ffffff",
   68584 => x"ffffff",
   68585 => x"ffffff",
   68586 => x"ffffff",
   68587 => x"ffffff",
   68588 => x"ffffff",
   68589 => x"ffffff",
   68590 => x"ffffff",
   68591 => x"ffffff",
   68592 => x"ffffff",
   68593 => x"ffffff",
   68594 => x"ffffff",
   68595 => x"ffffff",
   68596 => x"ffffff",
   68597 => x"ffffff",
   68598 => x"ffffff",
   68599 => x"ffffff",
   68600 => x"ffffff",
   68601 => x"ffffff",
   68602 => x"ffffff",
   68603 => x"ffffff",
   68604 => x"ffffff",
   68605 => x"ffffff",
   68606 => x"ffffff",
   68607 => x"ffffff",
   68608 => x"ffffff",
   68609 => x"ffffff",
   68610 => x"ffffff",
   68611 => x"ffffff",
   68612 => x"ffffff",
   68613 => x"ffffff",
   68614 => x"ffffff",
   68615 => x"ffffff",
   68616 => x"ffffff",
   68617 => x"ffffff",
   68618 => x"ffffff",
   68619 => x"ffffff",
   68620 => x"ffffff",
   68621 => x"ffffff",
   68622 => x"ffffff",
   68623 => x"ffffff",
   68624 => x"ffffff",
   68625 => x"ffffff",
   68626 => x"ffffff",
   68627 => x"ffffff",
   68628 => x"ffffff",
   68629 => x"ffffff",
   68630 => x"ffffff",
   68631 => x"ffffff",
   68632 => x"ffffff",
   68633 => x"ffffff",
   68634 => x"ffffff",
   68635 => x"ffffff",
   68636 => x"ffffff",
   68637 => x"ffffff",
   68638 => x"ffffff",
   68639 => x"ffffff",
   68640 => x"ffffff",
   68641 => x"ffffff",
   68642 => x"ffffff",
   68643 => x"ffffff",
   68644 => x"ffffff",
   68645 => x"ffffff",
   68646 => x"ffffff",
   68647 => x"ffffff",
   68648 => x"ffffff",
   68649 => x"ffffff",
   68650 => x"ffffff",
   68651 => x"ffffff",
   68652 => x"ffffff",
   68653 => x"ffffff",
   68654 => x"ffffff",
   68655 => x"ffffff",
   68656 => x"ffffff",
   68657 => x"ffffff",
   68658 => x"ffffff",
   68659 => x"ffffff",
   68660 => x"ffffff",
   68661 => x"ffffff",
   68662 => x"ffffff",
   68663 => x"ffffff",
   68664 => x"ffffff",
   68665 => x"ffffff",
   68666 => x"ffffff",
   68667 => x"ffffff",
   68668 => x"ffffff",
   68669 => x"ffffff",
   68670 => x"ffffff",
   68671 => x"ffffff",
   68672 => x"ffffff",
   68673 => x"ffffff",
   68674 => x"ffffff",
   68675 => x"ffffff",
   68676 => x"ffffff",
   68677 => x"ffffff",
   68678 => x"ffffff",
   68679 => x"ffffff",
   68680 => x"ffffff",
   68681 => x"ffffff",
   68682 => x"ffffff",
   68683 => x"ffffff",
   68684 => x"ffffff",
   68685 => x"ffffff",
   68686 => x"ffffff",
   68687 => x"ffffff",
   68688 => x"ffffff",
   68689 => x"ffffff",
   68690 => x"ffffff",
   68691 => x"ffffff",
   68692 => x"ffffff",
   68693 => x"ffffff",
   68694 => x"ffffff",
   68695 => x"ffffff",
   68696 => x"ffffff",
   68697 => x"ffffff",
   68698 => x"ffffff",
   68699 => x"ffffff",
   68700 => x"ffffff",
   68701 => x"ffffff",
   68702 => x"ffffff",
   68703 => x"ffffff",
   68704 => x"ffffff",
   68705 => x"ffffff",
   68706 => x"ffffff",
   68707 => x"ffffff",
   68708 => x"ffffff",
   68709 => x"ffffff",
   68710 => x"ffffff",
   68711 => x"ffffff",
   68712 => x"ffffff",
   68713 => x"ffffff",
   68714 => x"ffffff",
   68715 => x"ffffff",
   68716 => x"ffffff",
   68717 => x"ffffff",
   68718 => x"ffffff",
   68719 => x"ffffff",
   68720 => x"ffffff",
   68721 => x"ffffff",
   68722 => x"ffffff",
   68723 => x"ffffff",
   68724 => x"ffffff",
   68725 => x"ffffff",
   68726 => x"ffffff",
   68727 => x"ffffff",
   68728 => x"ffffff",
   68729 => x"ffffff",
   68730 => x"ffffff",
   68731 => x"ffffff",
   68732 => x"ffffff",
   68733 => x"ffffff",
   68734 => x"ffffff",
   68735 => x"ffffff",
   68736 => x"ffffff",
   68737 => x"ffffff",
   68738 => x"ffffff",
   68739 => x"ffffff",
   68740 => x"ffffff",
   68741 => x"ffffff",
   68742 => x"ffffff",
   68743 => x"ffffff",
   68744 => x"ffffff",
   68745 => x"ffffff",
   68746 => x"ffffff",
   68747 => x"ffffff",
   68748 => x"ffffff",
   68749 => x"ffffff",
   68750 => x"ffffff",
   68751 => x"ffffff",
   68752 => x"ffffff",
   68753 => x"ffffff",
   68754 => x"ffffff",
   68755 => x"ffffff",
   68756 => x"ffffff",
   68757 => x"ffffff",
   68758 => x"ffffff",
   68759 => x"ffffff",
   68760 => x"ffffff",
   68761 => x"ffffff",
   68762 => x"ffffff",
   68763 => x"ffffff",
   68764 => x"ffffff",
   68765 => x"ffffff",
   68766 => x"ffffff",
   68767 => x"ffffff",
   68768 => x"ffffff",
   68769 => x"ffffff",
   68770 => x"ffffff",
   68771 => x"ffffff",
   68772 => x"ffffff",
   68773 => x"ffffff",
   68774 => x"ffffff",
   68775 => x"ffffff",
   68776 => x"ffffff",
   68777 => x"ffffff",
   68778 => x"ffffff",
   68779 => x"ffffff",
   68780 => x"ffffff",
   68781 => x"ffffff",
   68782 => x"ffffff",
   68783 => x"ffffff",
   68784 => x"ffffff",
   68785 => x"ffffff",
   68786 => x"ffffff",
   68787 => x"ffffff",
   68788 => x"ffffff",
   68789 => x"ffffff",
   68790 => x"ffffff",
   68791 => x"ffffff",
   68792 => x"ffffff",
   68793 => x"ffffff",
   68794 => x"ffffff",
   68795 => x"ffffff",
   68796 => x"ffffff",
   68797 => x"ffffff",
   68798 => x"ffffff",
   68799 => x"ffffff",
   68800 => x"ffffff",
   68801 => x"ffffff",
   68802 => x"ffffff",
   68803 => x"ffffff",
   68804 => x"ffffff",
   68805 => x"ffffff",
   68806 => x"ffffff",
   68807 => x"ffffff",
   68808 => x"ffffff",
   68809 => x"ffffff",
   68810 => x"ffffff",
   68811 => x"ffffff",
   68812 => x"ffffff",
   68813 => x"ffffff",
   68814 => x"ffffff",
   68815 => x"ffffff",
   68816 => x"ffffff",
   68817 => x"ffffff",
   68818 => x"ffffff",
   68819 => x"ffffff",
   68820 => x"ffffff",
   68821 => x"ffffff",
   68822 => x"ffffff",
   68823 => x"ffffff",
   68824 => x"ffffff",
   68825 => x"ffffff",
   68826 => x"ffffff",
   68827 => x"ffffff",
   68828 => x"ffffff",
   68829 => x"ffffff",
   68830 => x"ffffff",
   68831 => x"ffffff",
   68832 => x"ffffff",
   68833 => x"ffffff",
   68834 => x"ffffff",
   68835 => x"ffffff",
   68836 => x"ffffff",
   68837 => x"ffffff",
   68838 => x"ffffff",
   68839 => x"ffffff",
   68840 => x"ffffff",
   68841 => x"ffffff",
   68842 => x"ffffff",
   68843 => x"ffffff",
   68844 => x"ffffff",
   68845 => x"ffffff",
   68846 => x"ffffff",
   68847 => x"ffffff",
   68848 => x"ffffff",
   68849 => x"ffffff",
   68850 => x"ffffff",
   68851 => x"ffffff",
   68852 => x"ffffff",
   68853 => x"ffffff",
   68854 => x"ffffff",
   68855 => x"ffffff",
   68856 => x"ffffff",
   68857 => x"ffffff",
   68858 => x"ffffff",
   68859 => x"ffffff",
   68860 => x"ffffff",
   68861 => x"ffffff",
   68862 => x"ffffff",
   68863 => x"ffffff",
   68864 => x"ffffff",
   68865 => x"ffffff",
   68866 => x"ffffff",
   68867 => x"ffffff",
   68868 => x"ffffff",
   68869 => x"ffffff",
   68870 => x"ffffff",
   68871 => x"ffffff",
   68872 => x"ffffff",
   68873 => x"ffffff",
   68874 => x"ffffff",
   68875 => x"ffffff",
   68876 => x"ffffff",
   68877 => x"ffffff",
   68878 => x"ffffff",
   68879 => x"ffffff",
   68880 => x"ffffff",
   68881 => x"ffffff",
   68882 => x"ffffff",
   68883 => x"ffffff",
   68884 => x"ffffff",
   68885 => x"ffffff",
   68886 => x"ffffff",
   68887 => x"ffffff",
   68888 => x"ffffff",
   68889 => x"ffffff",
   68890 => x"ffffff",
   68891 => x"ffffff",
   68892 => x"ffffff",
   68893 => x"ffffff",
   68894 => x"ffffff",
   68895 => x"ffffff",
   68896 => x"ffffff",
   68897 => x"ffffff",
   68898 => x"ffffff",
   68899 => x"ffffff",
   68900 => x"ffffff",
   68901 => x"ffffff",
   68902 => x"ffffff",
   68903 => x"ffffff",
   68904 => x"ffffff",
   68905 => x"ffffff",
   68906 => x"ffffff",
   68907 => x"ffffff",
   68908 => x"ffffff",
   68909 => x"ffffff",
   68910 => x"ffffff",
   68911 => x"ffffff",
   68912 => x"ffffff",
   68913 => x"ffffff",
   68914 => x"ffffff",
   68915 => x"ffffff",
   68916 => x"ffffff",
   68917 => x"ffffff",
   68918 => x"ffffff",
   68919 => x"ffffff",
   68920 => x"ffffff",
   68921 => x"ffffff",
   68922 => x"ffffff",
   68923 => x"ffffff",
   68924 => x"ffffff",
   68925 => x"ffffff",
   68926 => x"ffffff",
   68927 => x"ffffff",
   68928 => x"ffffff",
   68929 => x"ffffff",
   68930 => x"ffffff",
   68931 => x"ffffff",
   68932 => x"ffffff",
   68933 => x"ffffff",
   68934 => x"ffffff",
   68935 => x"ffffff",
   68936 => x"ffffff",
   68937 => x"ffffff",
   68938 => x"ffffff",
   68939 => x"ffffff",
   68940 => x"ffffff",
   68941 => x"ffffff",
   68942 => x"ffffff",
   68943 => x"ffffff",
   68944 => x"ffffff",
   68945 => x"ffffff",
   68946 => x"ffffff",
   68947 => x"ffffff",
   68948 => x"ffffff",
   68949 => x"ffffff",
   68950 => x"ffffff",
   68951 => x"ffffff",
   68952 => x"ffffff",
   68953 => x"ffffff",
   68954 => x"ffffff",
   68955 => x"ffffff",
   68956 => x"ffffff",
   68957 => x"ffffff",
   68958 => x"ffffff",
   68959 => x"ffffff",
   68960 => x"ffffff",
   68961 => x"ffffff",
   68962 => x"ffffff",
   68963 => x"ffffff",
   68964 => x"ffffff",
   68965 => x"ffffff",
   68966 => x"ffffff",
   68967 => x"ffffff",
   68968 => x"ffffff",
   68969 => x"ffffff",
   68970 => x"ffffff",
   68971 => x"ffffff",
   68972 => x"ffffff",
   68973 => x"ffffff",
   68974 => x"ffffff",
   68975 => x"ffffff",
   68976 => x"ffffff",
   68977 => x"ffffff",
   68978 => x"ffffff",
   68979 => x"ffffff",
   68980 => x"ffffff",
   68981 => x"ffffff",
   68982 => x"ffffff",
   68983 => x"ffffff",
   68984 => x"ffffff",
   68985 => x"ffffff",
   68986 => x"ffffff",
   68987 => x"ffffff",
   68988 => x"ffffff",
   68989 => x"ffffff",
   68990 => x"ffffff",
   68991 => x"ffffff",
   68992 => x"ffffff",
   68993 => x"ffffff",
   68994 => x"ffffff",
   68995 => x"ffffff",
   68996 => x"ffffff",
   68997 => x"ffffff",
   68998 => x"ffffff",
   68999 => x"ffffff",
   69000 => x"ffffff",
   69001 => x"ffffff",
   69002 => x"ffffff",
   69003 => x"ffffff",
   69004 => x"ffffff",
   69005 => x"ffffff",
   69006 => x"ffffff",
   69007 => x"ffffff",
   69008 => x"ffffff",
   69009 => x"ffffff",
   69010 => x"ffffff",
   69011 => x"ffffff",
   69012 => x"ffffff",
   69013 => x"ffffff",
   69014 => x"ffffff",
   69015 => x"ffffff",
   69016 => x"ffffff",
   69017 => x"ffffff",
   69018 => x"ffffff",
   69019 => x"ffffff",
   69020 => x"ffffff",
   69021 => x"ffffff",
   69022 => x"ffffff",
   69023 => x"ffffff",
   69024 => x"ffffff",
   69025 => x"ffffff",
   69026 => x"ffffff",
   69027 => x"ffffff",
   69028 => x"ffffff",
   69029 => x"ffffff",
   69030 => x"ffffff",
   69031 => x"ffffff",
   69032 => x"ffffff",
   69033 => x"ffffff",
   69034 => x"ffffff",
   69035 => x"ffffff",
   69036 => x"ffffff",
   69037 => x"ffffff",
   69038 => x"ffffff",
   69039 => x"ffffff",
   69040 => x"ffffff",
   69041 => x"ffffff",
   69042 => x"ffffff",
   69043 => x"ffffff",
   69044 => x"ffffff",
   69045 => x"ffffff",
   69046 => x"ffffff",
   69047 => x"ffffff",
   69048 => x"ffffff",
   69049 => x"ffffff",
   69050 => x"ffffff",
   69051 => x"ffffff",
   69052 => x"ffffff",
   69053 => x"ffffff",
   69054 => x"ffffff",
   69055 => x"ffffff",
   69056 => x"ffffff",
   69057 => x"ffffff",
   69058 => x"ffffff",
   69059 => x"ffffff",
   69060 => x"ffffff",
   69061 => x"ffffff",
   69062 => x"ffffff",
   69063 => x"ffffff",
   69064 => x"ffffff",
   69065 => x"ffffff",
   69066 => x"ffffff",
   69067 => x"ffffff",
   69068 => x"ffffff",
   69069 => x"ffffff",
   69070 => x"ffffff",
   69071 => x"ffffff",
   69072 => x"ffffff",
   69073 => x"ffffff",
   69074 => x"ffffff",
   69075 => x"ffffff",
   69076 => x"ffffff",
   69077 => x"ffffff",
   69078 => x"ffffff",
   69079 => x"ffffff",
   69080 => x"ffffff",
   69081 => x"ffffff",
   69082 => x"ffffff",
   69083 => x"ffffff",
   69084 => x"ffffff",
   69085 => x"ffffff",
   69086 => x"ffffff",
   69087 => x"ffffff",
   69088 => x"ffffff",
   69089 => x"ffffff",
   69090 => x"ffffff",
   69091 => x"ffffff",
   69092 => x"ffffff",
   69093 => x"ffffff",
   69094 => x"ffffff",
   69095 => x"ffffff",
   69096 => x"ffffff",
   69097 => x"ffffff",
   69098 => x"ffffff",
   69099 => x"ffffff",
   69100 => x"ffffff",
   69101 => x"ffffff",
   69102 => x"ffffff",
   69103 => x"ffffff",
   69104 => x"ffffff",
   69105 => x"ffffff",
   69106 => x"ffffff",
   69107 => x"ffffff",
   69108 => x"ffffff",
   69109 => x"ffffff",
   69110 => x"ffffff",
   69111 => x"ffffff",
   69112 => x"ffffff",
   69113 => x"ffffff",
   69114 => x"ffffff",
   69115 => x"ffffff",
   69116 => x"ffffff",
   69117 => x"ffffff",
   69118 => x"ffffff",
   69119 => x"ffffff",
   69120 => x"ffffff",
   69121 => x"ffffff",
   69122 => x"ffffff",
   69123 => x"ffffff",
   69124 => x"ffffff",
   69125 => x"ffffff",
   69126 => x"ffffff",
   69127 => x"ffffff",
   69128 => x"ffffff",
   69129 => x"ffffff",
   69130 => x"ffffff",
   69131 => x"ffffff",
   69132 => x"ffffff",
   69133 => x"ffffff",
   69134 => x"ffffff",
   69135 => x"ffffff",
   69136 => x"ffffff",
   69137 => x"ffffff",
   69138 => x"ffffff",
   69139 => x"ffffff",
   69140 => x"ffffff",
   69141 => x"ffffff",
   69142 => x"ffffff",
   69143 => x"ffffff",
   69144 => x"ffffff",
   69145 => x"ffffff",
   69146 => x"ffffff",
   69147 => x"ffffff",
   69148 => x"ffffff",
   69149 => x"ffffff",
   69150 => x"ffffff",
   69151 => x"ffffff",
   69152 => x"ffffff",
   69153 => x"ffffff",
   69154 => x"ffffff",
   69155 => x"ffffff",
   69156 => x"ffffff",
   69157 => x"ffffff",
   69158 => x"ffffff",
   69159 => x"ffffff",
   69160 => x"ffffff",
   69161 => x"ffffff",
   69162 => x"ffffff",
   69163 => x"ffffff",
   69164 => x"ffffff",
   69165 => x"ffffff",
   69166 => x"ffffff",
   69167 => x"ffffff",
   69168 => x"ffffff",
   69169 => x"ffffff",
   69170 => x"ffffff",
   69171 => x"ffffff",
   69172 => x"ffffff",
   69173 => x"ffffff",
   69174 => x"ffffff",
   69175 => x"ffffff",
   69176 => x"ffffff",
   69177 => x"ffffff",
   69178 => x"ffffff",
   69179 => x"ffffff",
   69180 => x"ffffff",
   69181 => x"ffffff",
   69182 => x"ffffff",
   69183 => x"ffffff",
   69184 => x"ffffff",
   69185 => x"ffffff",
   69186 => x"ffffff",
   69187 => x"ffffff",
   69188 => x"ffffff",
   69189 => x"ffffff",
   69190 => x"ffffff",
   69191 => x"ffffff",
   69192 => x"ffffff",
   69193 => x"ffffff",
   69194 => x"ffffff",
   69195 => x"ffffff",
   69196 => x"ffffff",
   69197 => x"ffffff",
   69198 => x"ffffff",
   69199 => x"ffffff",
   69200 => x"ffffff",
   69201 => x"ffffff",
   69202 => x"ffffff",
   69203 => x"ffffff",
   69204 => x"ffffff",
   69205 => x"ffffff",
   69206 => x"ffffff",
   69207 => x"ffffff",
   69208 => x"ffffff",
   69209 => x"ffffff",
   69210 => x"ffffff",
   69211 => x"ffffff",
   69212 => x"ffffff",
   69213 => x"ffffff",
   69214 => x"ffffff",
   69215 => x"ffffff",
   69216 => x"ffffff",
   69217 => x"ffffff",
   69218 => x"ffffff",
   69219 => x"ffffff",
   69220 => x"ffffff",
   69221 => x"ffffff",
   69222 => x"ffffff",
   69223 => x"ffffff",
   69224 => x"ffffff",
   69225 => x"ffffff",
   69226 => x"ffffff",
   69227 => x"ffffff",
   69228 => x"ffffff",
   69229 => x"ffffff",
   69230 => x"ffffff",
   69231 => x"ffffff",
   69232 => x"ffffff",
   69233 => x"ffffff",
   69234 => x"ffffff",
   69235 => x"ffffff",
   69236 => x"ffffff",
   69237 => x"ffffff",
   69238 => x"ffffff",
   69239 => x"ffffff",
   69240 => x"ffffff",
   69241 => x"ffffff",
   69242 => x"ffffff",
   69243 => x"ffffff",
   69244 => x"ffffff",
   69245 => x"ffffff",
   69246 => x"ffffff",
   69247 => x"ffffff",
   69248 => x"ffffff",
   69249 => x"ffffff",
   69250 => x"ffffff",
   69251 => x"ffffff",
   69252 => x"ffffff",
   69253 => x"ffffff",
   69254 => x"ffffff",
   69255 => x"ffffff",
   69256 => x"ffffff",
   69257 => x"ffffff",
   69258 => x"ffffff",
   69259 => x"ffffff",
   69260 => x"ffffff",
   69261 => x"ffffff",
   69262 => x"ffffff",
   69263 => x"ffffff",
   69264 => x"ffffff",
   69265 => x"ffffff",
   69266 => x"ffffff",
   69267 => x"ffffff",
   69268 => x"ffffff",
   69269 => x"ffffff",
   69270 => x"ffffff",
   69271 => x"ffffff",
   69272 => x"ffffff",
   69273 => x"ffffff",
   69274 => x"ffffff",
   69275 => x"ffffff",
   69276 => x"ffffff",
   69277 => x"ffffff",
   69278 => x"ffffff",
   69279 => x"ffffff",
   69280 => x"ffffff",
   69281 => x"ffffff",
   69282 => x"ffffff",
   69283 => x"ffffff",
   69284 => x"ffffff",
   69285 => x"ffffff",
   69286 => x"ffffff",
   69287 => x"ffffff",
   69288 => x"ffffff",
   69289 => x"ffffff",
   69290 => x"ffffff",
   69291 => x"ffffff",
   69292 => x"ffffff",
   69293 => x"ffffff",
   69294 => x"ffffff",
   69295 => x"ffffff",
   69296 => x"ffffff",
   69297 => x"ffffff",
   69298 => x"ffffff",
   69299 => x"ffffff",
   69300 => x"ffffff",
   69301 => x"ffffff",
   69302 => x"ffffff",
   69303 => x"ffffff",
   69304 => x"ffffff",
   69305 => x"ffffff",
   69306 => x"ffffff",
   69307 => x"ffffff",
   69308 => x"ffffff",
   69309 => x"ffffff",
   69310 => x"ffffff",
   69311 => x"ffffff",
   69312 => x"ffffff",
   69313 => x"ffffff",
   69314 => x"ffffff",
   69315 => x"ffffff",
   69316 => x"ffffff",
   69317 => x"ffffff",
   69318 => x"ffffff",
   69319 => x"ffffff",
   69320 => x"ffffff",
   69321 => x"ffffff",
   69322 => x"ffffff",
   69323 => x"ffffff",
   69324 => x"ffffff",
   69325 => x"ffffff",
   69326 => x"ffffff",
   69327 => x"ffffff",
   69328 => x"ffffff",
   69329 => x"ffffff",
   69330 => x"ffffff",
   69331 => x"ffffff",
   69332 => x"ffffff",
   69333 => x"ffffff",
   69334 => x"ffffff",
   69335 => x"ffffff",
   69336 => x"ffffff",
   69337 => x"ffffff",
   69338 => x"ffffff",
   69339 => x"ffffff",
   69340 => x"ffffff",
   69341 => x"ffffff",
   69342 => x"ffffff",
   69343 => x"ffffff",
   69344 => x"ffffff",
   69345 => x"ffffff",
   69346 => x"ffffff",
   69347 => x"ffffff",
   69348 => x"ffffff",
   69349 => x"ffffff",
   69350 => x"ffffff",
   69351 => x"ffffff",
   69352 => x"ffffff",
   69353 => x"ffffff",
   69354 => x"ffffff",
   69355 => x"ffffff",
   69356 => x"ffffff",
   69357 => x"ffffff",
   69358 => x"ffffff",
   69359 => x"ffffff",
   69360 => x"ffffff",
   69361 => x"ffffff",
   69362 => x"ffffff",
   69363 => x"ffffff",
   69364 => x"ffffff",
   69365 => x"ffffff",
   69366 => x"ffffff",
   69367 => x"ffffff",
   69368 => x"ffffff",
   69369 => x"ffffff",
   69370 => x"ffffff",
   69371 => x"ffffff",
   69372 => x"ffffff",
   69373 => x"ffffff",
   69374 => x"ffffff",
   69375 => x"ffffff",
   69376 => x"ffffff",
   69377 => x"ffffff",
   69378 => x"ffffff",
   69379 => x"ffffff",
   69380 => x"ffffff",
   69381 => x"ffffff",
   69382 => x"ffffff",
   69383 => x"ffffff",
   69384 => x"ffffff",
   69385 => x"ffffff",
   69386 => x"ffffff",
   69387 => x"ffffff",
   69388 => x"ffffff",
   69389 => x"ffffff",
   69390 => x"ffffff",
   69391 => x"ffffff",
   69392 => x"ffffff",
   69393 => x"ffffff",
   69394 => x"ffffff",
   69395 => x"ffffff",
   69396 => x"ffffff",
   69397 => x"ffffff",
   69398 => x"ffffff",
   69399 => x"ffffff",
   69400 => x"ffffff",
   69401 => x"ffffff",
   69402 => x"ffffff",
   69403 => x"ffffff",
   69404 => x"ffffff",
   69405 => x"ffffff",
   69406 => x"ffffff",
   69407 => x"ffffff",
   69408 => x"ffffff",
   69409 => x"ffffff",
   69410 => x"ffffff",
   69411 => x"ffffff",
   69412 => x"ffffff",
   69413 => x"ffffff",
   69414 => x"ffffff",
   69415 => x"ffffff",
   69416 => x"ffffff",
   69417 => x"ffffff",
   69418 => x"ffffff",
   69419 => x"ffffff",
   69420 => x"ffffff",
   69421 => x"ffffff",
   69422 => x"ffffff",
   69423 => x"ffffff",
   69424 => x"ffffff",
   69425 => x"ffffff",
   69426 => x"ffffff",
   69427 => x"ffffff",
   69428 => x"ffffff",
   69429 => x"ffffff",
   69430 => x"ffffff",
   69431 => x"ffffff",
   69432 => x"ffffff",
   69433 => x"ffffff",
   69434 => x"ffffff",
   69435 => x"ffffff",
   69436 => x"ffffff",
   69437 => x"ffffff",
   69438 => x"ffffff",
   69439 => x"ffffff",
   69440 => x"ffffff",
   69441 => x"ffffff",
   69442 => x"ffffff",
   69443 => x"ffffff",
   69444 => x"ffffff",
   69445 => x"ffffff",
   69446 => x"ffffff",
   69447 => x"ffffff",
   69448 => x"ffffff",
   69449 => x"ffffff",
   69450 => x"ffffff",
   69451 => x"ffffff",
   69452 => x"ffffff",
   69453 => x"ffffff",
   69454 => x"ffffff",
   69455 => x"ffffff",
   69456 => x"ffffff",
   69457 => x"ffffff",
   69458 => x"ffffff",
   69459 => x"ffffff",
   69460 => x"ffffff",
   69461 => x"ffffff",
   69462 => x"ffffff",
   69463 => x"ffffff",
   69464 => x"ffffff",
   69465 => x"ffffff",
   69466 => x"ffffff",
   69467 => x"ffffff",
   69468 => x"ffffff",
   69469 => x"ffffff",
   69470 => x"ffffff",
   69471 => x"ffffff",
   69472 => x"ffffff",
   69473 => x"ffffff",
   69474 => x"ffffff",
   69475 => x"ffffff",
   69476 => x"ffffff",
   69477 => x"ffffff",
   69478 => x"ffffff",
   69479 => x"ffffff",
   69480 => x"ffffff",
   69481 => x"ffffff",
   69482 => x"ffffff",
   69483 => x"ffffff",
   69484 => x"ffffff",
   69485 => x"ffffff",
   69486 => x"ffffff",
   69487 => x"ffffff",
   69488 => x"ffffff",
   69489 => x"ffffff",
   69490 => x"ffffff",
   69491 => x"ffffff",
   69492 => x"ffffff",
   69493 => x"ffffff",
   69494 => x"ffffff",
   69495 => x"ffffff",
   69496 => x"ffffff",
   69497 => x"ffffff",
   69498 => x"ffffff",
   69499 => x"ffffff",
   69500 => x"ffffff",
   69501 => x"ffffff",
   69502 => x"ffffff",
   69503 => x"ffffff",
   69504 => x"ffffff",
   69505 => x"ffffff",
   69506 => x"ffffff",
   69507 => x"ffffff",
   69508 => x"ffffff",
   69509 => x"ffffff",
   69510 => x"ffffff",
   69511 => x"ffffff",
   69512 => x"ffffff",
   69513 => x"ffffff",
   69514 => x"ffffff",
   69515 => x"ffffff",
   69516 => x"ffffff",
   69517 => x"ffffff",
   69518 => x"ffffff",
   69519 => x"ffffff",
   69520 => x"ffffff",
   69521 => x"ffffff",
   69522 => x"ffffff",
   69523 => x"ffffff",
   69524 => x"ffffff",
   69525 => x"ffffff",
   69526 => x"ffffff",
   69527 => x"ffffff",
   69528 => x"ffffff",
   69529 => x"ffffff",
   69530 => x"ffffff",
   69531 => x"ffffff",
   69532 => x"ffffff",
   69533 => x"ffffff",
   69534 => x"ffffff",
   69535 => x"ffffff",
   69536 => x"ffffff",
   69537 => x"ffffff",
   69538 => x"ffffff",
   69539 => x"ffffff",
   69540 => x"ffffff",
   69541 => x"ffffff",
   69542 => x"ffffff",
   69543 => x"ffffff",
   69544 => x"ffffff",
   69545 => x"ffffff",
   69546 => x"ffffff",
   69547 => x"ffffff",
   69548 => x"ffffff",
   69549 => x"ffffff",
   69550 => x"ffffff",
   69551 => x"ffffff",
   69552 => x"ffffff",
   69553 => x"ffffff",
   69554 => x"ffffff",
   69555 => x"ffffff",
   69556 => x"ffffff",
   69557 => x"ffffff",
   69558 => x"ffffff",
   69559 => x"ffffff",
   69560 => x"ffffff",
   69561 => x"ffffff",
   69562 => x"ffffff",
   69563 => x"ffffff",
   69564 => x"ffffff",
   69565 => x"ffffff",
   69566 => x"ffffff",
   69567 => x"ffffff",
   69568 => x"ffffff",
   69569 => x"ffffff",
   69570 => x"ffffff",
   69571 => x"ffffff",
   69572 => x"ffffff",
   69573 => x"ffffff",
   69574 => x"ffffff",
   69575 => x"ffffff",
   69576 => x"ffffff",
   69577 => x"ffffff",
   69578 => x"ffffff",
   69579 => x"ffffff",
   69580 => x"ffffff",
   69581 => x"ffffff",
   69582 => x"ffffff",
   69583 => x"ffffff",
   69584 => x"ffffff",
   69585 => x"ffffff",
   69586 => x"ffffff",
   69587 => x"ffffff",
   69588 => x"ffffff",
   69589 => x"ffffff",
   69590 => x"ffffff",
   69591 => x"ffffff",
   69592 => x"ffffff",
   69593 => x"ffffff",
   69594 => x"ffffff",
   69595 => x"ffffff",
   69596 => x"ffffff",
   69597 => x"ffffff",
   69598 => x"ffffff",
   69599 => x"ffffff",
   69600 => x"ffffff",
   69601 => x"ffffff",
   69602 => x"ffffff",
   69603 => x"ffffff",
   69604 => x"ffffff",
   69605 => x"ffffff",
   69606 => x"ffffff",
   69607 => x"ffffff",
   69608 => x"ffffff",
   69609 => x"ffffff",
   69610 => x"ffffff",
   69611 => x"ffffff",
   69612 => x"ffffff",
   69613 => x"ffffff",
   69614 => x"ffffff",
   69615 => x"ffffff",
   69616 => x"ffffff",
   69617 => x"ffffff",
   69618 => x"ffffff",
   69619 => x"ffffff",
   69620 => x"ffffff",
   69621 => x"ffffff",
   69622 => x"ffffff",
   69623 => x"ffffff",
   69624 => x"ffffff",
   69625 => x"ffffff",
   69626 => x"ffffff",
   69627 => x"ffffff",
   69628 => x"ffffff",
   69629 => x"ffffff",
   69630 => x"ffffff",
   69631 => x"ffffff",
   69632 => x"ffffff",
   69633 => x"ffffff",
   69634 => x"ffffff",
   69635 => x"ffffff",
   69636 => x"ffffff",
   69637 => x"ffffff",
   69638 => x"ffffff",
   69639 => x"ffffff",
   69640 => x"ffffff",
   69641 => x"ffffff",
   69642 => x"ffffff",
   69643 => x"ffffff",
   69644 => x"ffffff",
   69645 => x"ffffff",
   69646 => x"ffffff",
   69647 => x"ffffff",
   69648 => x"ffffff",
   69649 => x"ffffff",
   69650 => x"ffffff",
   69651 => x"ffffff",
   69652 => x"ffffff",
   69653 => x"ffffff",
   69654 => x"ffffff",
   69655 => x"ffffff",
   69656 => x"ffffff",
   69657 => x"ffffff",
   69658 => x"ffffff",
   69659 => x"ffffff",
   69660 => x"ffffff",
   69661 => x"ffffff",
   69662 => x"ffffff",
   69663 => x"ffffff",
   69664 => x"ffffff",
   69665 => x"ffffff",
   69666 => x"ffffff",
   69667 => x"ffffff",
   69668 => x"ffffff",
   69669 => x"ffffff",
   69670 => x"ffffff",
   69671 => x"ffffff",
   69672 => x"ffffff",
   69673 => x"ffffff",
   69674 => x"ffffff",
   69675 => x"ffffff",
   69676 => x"ffffff",
   69677 => x"ffffff",
   69678 => x"ffffff",
   69679 => x"ffffff",
   69680 => x"ffffff",
   69681 => x"ffffff",
   69682 => x"ffffff",
   69683 => x"ffffff",
   69684 => x"ffffff",
   69685 => x"ffffff",
   69686 => x"ffffff",
   69687 => x"ffffff",
   69688 => x"ffffff",
   69689 => x"ffffff",
   69690 => x"ffffff",
   69691 => x"ffffff",
   69692 => x"ffffff",
   69693 => x"ffffff",
   69694 => x"ffffff",
   69695 => x"ffffff",
   69696 => x"ffffff",
   69697 => x"ffffff",
   69698 => x"ffffff",
   69699 => x"ffffff",
   69700 => x"ffffff",
   69701 => x"ffffff",
   69702 => x"ffffff",
   69703 => x"ffffff",
   69704 => x"ffffff",
   69705 => x"ffffff",
   69706 => x"ffffff",
   69707 => x"ffffff",
   69708 => x"ffffff",
   69709 => x"ffffff",
   69710 => x"ffffff",
   69711 => x"ffffff",
   69712 => x"ffffff",
   69713 => x"ffffff",
   69714 => x"ffffff",
   69715 => x"ffffff",
   69716 => x"ffffff",
   69717 => x"ffffff",
   69718 => x"ffffff",
   69719 => x"ffffff",
   69720 => x"ffffff",
   69721 => x"ffffff",
   69722 => x"ffffff",
   69723 => x"ffffff",
   69724 => x"ffffff",
   69725 => x"ffffff",
   69726 => x"ffffff",
   69727 => x"ffffff",
   69728 => x"ffffff",
   69729 => x"ffffff",
   69730 => x"ffffff",
   69731 => x"ffffff",
   69732 => x"ffffff",
   69733 => x"ffffff",
   69734 => x"ffffff",
   69735 => x"ffffff",
   69736 => x"ffffff",
   69737 => x"ffffff",
   69738 => x"ffffff",
   69739 => x"ffffff",
   69740 => x"ffffff",
   69741 => x"ffffff",
   69742 => x"ffffff",
   69743 => x"ffffff",
   69744 => x"ffffff",
   69745 => x"ffffff",
   69746 => x"ffffff",
   69747 => x"ffffff",
   69748 => x"ffffff",
   69749 => x"ffffff",
   69750 => x"ffffff",
   69751 => x"ffffff",
   69752 => x"ffffff",
   69753 => x"ffffff",
   69754 => x"ffffff",
   69755 => x"ffffff",
   69756 => x"ffffff",
   69757 => x"ffffff",
   69758 => x"ffffff",
   69759 => x"ffffff",
   69760 => x"ffffff",
   69761 => x"ffffff",
   69762 => x"ffffff",
   69763 => x"ffffff",
   69764 => x"ffffff",
   69765 => x"ffffff",
   69766 => x"ffffff",
   69767 => x"ffffff",
   69768 => x"ffffff",
   69769 => x"ffffff",
   69770 => x"ffffff",
   69771 => x"ffffff",
   69772 => x"ffffff",
   69773 => x"ffffff",
   69774 => x"ffffff",
   69775 => x"ffffff",
   69776 => x"ffffff",
   69777 => x"ffffff",
   69778 => x"ffffff",
   69779 => x"ffffff",
   69780 => x"ffffff",
   69781 => x"ffffff",
   69782 => x"ffffff",
   69783 => x"ffffff",
   69784 => x"ffffff",
   69785 => x"ffffff",
   69786 => x"ffffff",
   69787 => x"ffffff",
   69788 => x"ffffff",
   69789 => x"ffffff",
   69790 => x"ffffff",
   69791 => x"ffffff",
   69792 => x"ffffff",
   69793 => x"ffffff",
   69794 => x"ffffff",
   69795 => x"ffffff",
   69796 => x"ffffff",
   69797 => x"ffffff",
   69798 => x"ffffff",
   69799 => x"ffffff",
   69800 => x"ffffff",
   69801 => x"ffffff",
   69802 => x"ffffff",
   69803 => x"ffffff",
   69804 => x"ffffff",
   69805 => x"ffffff",
   69806 => x"ffffff",
   69807 => x"ffffff",
   69808 => x"ffffff",
   69809 => x"ffffff",
   69810 => x"ffffff",
   69811 => x"ffffff",
   69812 => x"ffffff",
   69813 => x"ffffff",
   69814 => x"ffffff",
   69815 => x"ffffff",
   69816 => x"ffffff",
   69817 => x"ffffff",
   69818 => x"ffffff",
   69819 => x"ffffff",
   69820 => x"ffffff",
   69821 => x"ffffff",
   69822 => x"ffffff",
   69823 => x"ffffff",
   69824 => x"ffffff",
   69825 => x"ffffff",
   69826 => x"ffffff",
   69827 => x"ffffff",
   69828 => x"ffffff",
   69829 => x"ffffff",
   69830 => x"ffffff",
   69831 => x"ffffff",
   69832 => x"ffffff",
   69833 => x"ffffff",
   69834 => x"ffffff",
   69835 => x"ffffff",
   69836 => x"ffffff",
   69837 => x"ffffff",
   69838 => x"ffffff",
   69839 => x"ffffff",
   69840 => x"ffffff",
   69841 => x"ffffff",
   69842 => x"ffffff",
   69843 => x"ffffff",
   69844 => x"ffffff",
   69845 => x"ffffff",
   69846 => x"ffffff",
   69847 => x"ffffff",
   69848 => x"ffffff",
   69849 => x"ffffff",
   69850 => x"ffffff",
   69851 => x"ffffff",
   69852 => x"ffffff",
   69853 => x"ffffff",
   69854 => x"ffffff",
   69855 => x"ffffff",
   69856 => x"ffffff",
   69857 => x"ffffff",
   69858 => x"ffffff",
   69859 => x"ffffff",
   69860 => x"ffffff",
   69861 => x"ffffff",
   69862 => x"ffffff",
   69863 => x"ffffff",
   69864 => x"ffffff",
   69865 => x"ffffff",
   69866 => x"ffffff",
   69867 => x"ffffff",
   69868 => x"ffffff",
   69869 => x"ffffff",
   69870 => x"ffffff",
   69871 => x"ffffff",
   69872 => x"ffffff",
   69873 => x"ffffff",
   69874 => x"ffffff",
   69875 => x"ffffff",
   69876 => x"ffffff",
   69877 => x"ffffff",
   69878 => x"ffffff",
   69879 => x"ffffff",
   69880 => x"ffffff",
   69881 => x"ffffff",
   69882 => x"ffffff",
   69883 => x"ffffff",
   69884 => x"ffffff",
   69885 => x"ffffff",
   69886 => x"ffffff",
   69887 => x"ffffff",
   69888 => x"ffffff",
   69889 => x"ffffff",
   69890 => x"ffffff",
   69891 => x"ffffff",
   69892 => x"ffffff",
   69893 => x"ffffff",
   69894 => x"ffffff",
   69895 => x"ffffff",
   69896 => x"ffffff",
   69897 => x"ffffff",
   69898 => x"ffffff",
   69899 => x"ffffff",
   69900 => x"ffffff",
   69901 => x"ffffff",
   69902 => x"ffffff",
   69903 => x"ffffff",
   69904 => x"ffffff",
   69905 => x"ffffff",
   69906 => x"ffffff",
   69907 => x"ffffff",
   69908 => x"ffffff",
   69909 => x"ffffff",
   69910 => x"ffffff",
   69911 => x"ffffff",
   69912 => x"ffffff",
   69913 => x"ffffff",
   69914 => x"ffffff",
   69915 => x"ffffff",
   69916 => x"ffffff",
   69917 => x"ffffff",
   69918 => x"ffffff",
   69919 => x"ffffff",
   69920 => x"ffffff",
   69921 => x"ffffff",
   69922 => x"ffffff",
   69923 => x"ffffff",
   69924 => x"ffffff",
   69925 => x"ffffff",
   69926 => x"ffffff",
   69927 => x"ffffff",
   69928 => x"ffffff",
   69929 => x"ffffff",
   69930 => x"ffffff",
   69931 => x"ffffff",
   69932 => x"ffffff",
   69933 => x"ffffff",
   69934 => x"ffffff",
   69935 => x"ffffff",
   69936 => x"ffffff",
   69937 => x"ffffff",
   69938 => x"ffffff",
   69939 => x"ffffff",
   69940 => x"ffffff",
   69941 => x"ffffff",
   69942 => x"ffffff",
   69943 => x"ffffff",
   69944 => x"ffffff",
   69945 => x"ffffff",
   69946 => x"ffffff",
   69947 => x"ffffff",
   69948 => x"ffffff",
   69949 => x"ffffff",
   69950 => x"ffffff",
   69951 => x"ffffff",
   69952 => x"ffffff",
   69953 => x"ffffff",
   69954 => x"ffffff",
   69955 => x"ffffff",
   69956 => x"ffffff",
   69957 => x"ffffff",
   69958 => x"ffffff",
   69959 => x"ffffff",
   69960 => x"ffffff",
   69961 => x"ffffff",
   69962 => x"ffffff",
   69963 => x"ffffff",
   69964 => x"ffffff",
   69965 => x"ffffff",
   69966 => x"ffffff",
   69967 => x"ffffff",
   69968 => x"ffffff",
   69969 => x"ffffff",
   69970 => x"ffffff",
   69971 => x"ffffff",
   69972 => x"ffffff",
   69973 => x"ffffff",
   69974 => x"ffffff",
   69975 => x"ffffff",
   69976 => x"ffffff",
   69977 => x"ffffff",
   69978 => x"ffffff",
   69979 => x"ffffff",
   69980 => x"ffffff",
   69981 => x"ffffff",
   69982 => x"ffffff",
   69983 => x"ffffff",
   69984 => x"ffffff",
   69985 => x"ffffff",
   69986 => x"ffffff",
   69987 => x"ffffff",
   69988 => x"ffffff",
   69989 => x"ffffff",
   69990 => x"ffffff",
   69991 => x"ffffff",
   69992 => x"ffffff",
   69993 => x"ffffff",
   69994 => x"ffffff",
   69995 => x"ffffff",
   69996 => x"ffffff",
   69997 => x"ffffff",
   69998 => x"ffffff",
   69999 => x"ffffff",
   70000 => x"ffffff",
   70001 => x"ffffff",
   70002 => x"ffffff",
   70003 => x"ffffff",
   70004 => x"ffffff",
   70005 => x"ffffff",
   70006 => x"ffffff",
   70007 => x"ffffff",
   70008 => x"ffffff",
   70009 => x"ffffff",
   70010 => x"ffffff",
   70011 => x"ffffff",
   70012 => x"ffffff",
   70013 => x"ffffff",
   70014 => x"ffffff",
   70015 => x"ffffff",
   70016 => x"ffffff",
   70017 => x"ffffff",
   70018 => x"ffffff",
   70019 => x"ffffff",
   70020 => x"ffffff",
   70021 => x"ffffff",
   70022 => x"ffffff",
   70023 => x"ffffff",
   70024 => x"ffffff",
   70025 => x"ffffff",
   70026 => x"ffffff",
   70027 => x"ffffff",
   70028 => x"ffffff",
   70029 => x"ffffff",
   70030 => x"ffffff",
   70031 => x"ffffff",
   70032 => x"ffffff",
   70033 => x"ffffff",
   70034 => x"ffffff",
   70035 => x"ffffff",
   70036 => x"ffffff",
   70037 => x"ffffff",
   70038 => x"ffffff",
   70039 => x"ffffff",
   70040 => x"ffffff",
   70041 => x"ffffff",
   70042 => x"ffffff",
   70043 => x"ffffff",
   70044 => x"ffffff",
   70045 => x"ffffff",
   70046 => x"ffffff",
   70047 => x"ffffff",
   70048 => x"ffffff",
   70049 => x"ffffff",
   70050 => x"ffffff",
   70051 => x"ffffff",
   70052 => x"ffffff",
   70053 => x"ffffff",
   70054 => x"ffffff",
   70055 => x"ffffff",
   70056 => x"ffffff",
   70057 => x"ffffff",
   70058 => x"ffffff",
   70059 => x"ffffff",
   70060 => x"ffffff",
   70061 => x"ffffff",
   70062 => x"ffffff",
   70063 => x"ffffff",
   70064 => x"ffffff",
   70065 => x"ffffff",
   70066 => x"ffffff",
   70067 => x"ffffff",
   70068 => x"ffffff",
   70069 => x"ffffff",
   70070 => x"ffffff",
   70071 => x"ffffff",
   70072 => x"ffffff",
   70073 => x"ffffff",
   70074 => x"ffffff",
   70075 => x"ffffff",
   70076 => x"ffffff",
   70077 => x"ffffff",
   70078 => x"ffffff",
   70079 => x"ffffff",
   70080 => x"ffffff",
   70081 => x"ffffff",
   70082 => x"ffffff",
   70083 => x"ffffff",
   70084 => x"ffffff",
   70085 => x"ffffff",
   70086 => x"ffffff",
   70087 => x"ffffff",
   70088 => x"ffffff",
   70089 => x"ffffff",
   70090 => x"ffffff",
   70091 => x"ffffff",
   70092 => x"ffffff",
   70093 => x"ffffff",
   70094 => x"ffffff",
   70095 => x"ffffff",
   70096 => x"ffffff",
   70097 => x"ffffff",
   70098 => x"ffffff",
   70099 => x"ffffff",
   70100 => x"ffffff",
   70101 => x"ffffff",
   70102 => x"ffffff",
   70103 => x"ffffff",
   70104 => x"ffffff",
   70105 => x"ffffff",
   70106 => x"ffffff",
   70107 => x"ffffff",
   70108 => x"ffffff",
   70109 => x"ffffff",
   70110 => x"ffffff",
   70111 => x"ffffff",
   70112 => x"ffffff",
   70113 => x"ffffff",
   70114 => x"ffffff",
   70115 => x"ffffff",
   70116 => x"ffffff",
   70117 => x"ffffff",
   70118 => x"ffffff",
   70119 => x"ffffff",
   70120 => x"ffffff",
   70121 => x"ffffff",
   70122 => x"ffffff",
   70123 => x"ffffff",
   70124 => x"ffffff",
   70125 => x"ffffff",
   70126 => x"ffffff",
   70127 => x"ffffff",
   70128 => x"ffffff",
   70129 => x"ffffff",
   70130 => x"ffffff",
   70131 => x"ffffff",
   70132 => x"ffffff",
   70133 => x"ffffff",
   70134 => x"ffffff",
   70135 => x"ffffff",
   70136 => x"ffffff",
   70137 => x"ffffff",
   70138 => x"ffffff",
   70139 => x"ffffff",
   70140 => x"ffffff",
   70141 => x"ffffff",
   70142 => x"ffffff",
   70143 => x"ffffff",
   70144 => x"ffffff",
   70145 => x"ffffff",
   70146 => x"ffffff",
   70147 => x"ffffff",
   70148 => x"ffffff",
   70149 => x"ffffff",
   70150 => x"ffffff",
   70151 => x"ffffff",
   70152 => x"ffffff",
   70153 => x"ffffff",
   70154 => x"ffffff",
   70155 => x"ffffff",
   70156 => x"ffffff",
   70157 => x"ffffff",
   70158 => x"ffffff",
   70159 => x"ffffff",
   70160 => x"ffffff",
   70161 => x"ffffff",
   70162 => x"ffffff",
   70163 => x"ffffff",
   70164 => x"ffffff",
   70165 => x"ffffff",
   70166 => x"ffffff",
   70167 => x"ffffff",
   70168 => x"ffffff",
   70169 => x"ffffff",
   70170 => x"ffffff",
   70171 => x"ffffff",
   70172 => x"ffffff",
   70173 => x"ffffff",
   70174 => x"ffffff",
   70175 => x"ffffff",
   70176 => x"ffffff",
   70177 => x"ffffff",
   70178 => x"ffffff",
   70179 => x"ffffff",
   70180 => x"ffffff",
   70181 => x"ffffff",
   70182 => x"ffffff",
   70183 => x"ffffff",
   70184 => x"ffffff",
   70185 => x"ffffff",
   70186 => x"ffffff",
   70187 => x"ffffff",
   70188 => x"ffffff",
   70189 => x"ffffff",
   70190 => x"ffffff",
   70191 => x"ffffff",
   70192 => x"ffffff",
   70193 => x"ffffff",
   70194 => x"ffffff",
   70195 => x"ffffff",
   70196 => x"ffffff",
   70197 => x"ffffff",
   70198 => x"ffffff",
   70199 => x"ffffff",
   70200 => x"ffffff",
   70201 => x"ffffff",
   70202 => x"ffffff",
   70203 => x"ffffff",
   70204 => x"ffffff",
   70205 => x"ffffff",
   70206 => x"ffffff",
   70207 => x"ffffff",
   70208 => x"ffffff",
   70209 => x"ffffff",
   70210 => x"ffffff",
   70211 => x"ffffff",
   70212 => x"ffffff",
   70213 => x"ffffff",
   70214 => x"ffffff",
   70215 => x"ffffff",
   70216 => x"ffffff",
   70217 => x"ffffff",
   70218 => x"ffffff",
   70219 => x"ffffff",
   70220 => x"ffffff",
   70221 => x"ffffff",
   70222 => x"ffffff",
   70223 => x"ffffff",
   70224 => x"ffffff",
   70225 => x"ffffff",
   70226 => x"ffffff",
   70227 => x"ffffff",
   70228 => x"ffffff",
   70229 => x"ffffff",
   70230 => x"ffffff",
   70231 => x"ffffff",
   70232 => x"ffffff",
   70233 => x"ffffff",
   70234 => x"ffffff",
   70235 => x"ffffff",
   70236 => x"ffffff",
   70237 => x"ffffff",
   70238 => x"ffffff",
   70239 => x"ffffff",
   70240 => x"ffffff",
   70241 => x"ffffff",
   70242 => x"ffffff",
   70243 => x"ffffff",
   70244 => x"ffffff",
   70245 => x"ffffff",
   70246 => x"ffffff",
   70247 => x"ffffff",
   70248 => x"ffffff",
   70249 => x"ffffff",
   70250 => x"ffffff",
   70251 => x"ffffff",
   70252 => x"ffffff",
   70253 => x"ffffff",
   70254 => x"ffffff",
   70255 => x"ffffff",
   70256 => x"ffffff",
   70257 => x"ffffff",
   70258 => x"ffffff",
   70259 => x"ffffff",
   70260 => x"ffffff",
   70261 => x"ffffff",
   70262 => x"ffffff",
   70263 => x"ffffff",
   70264 => x"ffffff",
   70265 => x"ffffff",
   70266 => x"ffffff",
   70267 => x"ffffff",
   70268 => x"ffffff",
   70269 => x"ffffff",
   70270 => x"ffffff",
   70271 => x"ffffff",
   70272 => x"ffffff",
   70273 => x"ffffff",
   70274 => x"ffffff",
   70275 => x"ffffff",
   70276 => x"ffffff",
   70277 => x"ffffff",
   70278 => x"ffffff",
   70279 => x"ffffff",
   70280 => x"ffffff",
   70281 => x"ffffff",
   70282 => x"ffffff",
   70283 => x"ffffff",
   70284 => x"ffffff",
   70285 => x"ffffff",
   70286 => x"ffffff",
   70287 => x"ffffff",
   70288 => x"ffffff",
   70289 => x"ffffff",
   70290 => x"ffffff",
   70291 => x"ffffff",
   70292 => x"ffffff",
   70293 => x"ffffff",
   70294 => x"ffffff",
   70295 => x"ffffff",
   70296 => x"ffffff",
   70297 => x"ffffff",
   70298 => x"ffffff",
   70299 => x"ffffff",
   70300 => x"ffffff",
   70301 => x"ffffff",
   70302 => x"ffffff",
   70303 => x"ffffff",
   70304 => x"ffffff",
   70305 => x"ffffff",
   70306 => x"ffffff",
   70307 => x"ffffff",
   70308 => x"ffffff",
   70309 => x"ffffff",
   70310 => x"ffffff",
   70311 => x"ffffff",
   70312 => x"ffffff",
   70313 => x"ffffff",
   70314 => x"ffffff",
   70315 => x"ffffff",
   70316 => x"ffffff",
   70317 => x"ffffff",
   70318 => x"ffffff",
   70319 => x"ffffff",
   70320 => x"ffffff",
   70321 => x"ffffff",
   70322 => x"ffffff",
   70323 => x"ffffff",
   70324 => x"ffffff",
   70325 => x"ffffff",
   70326 => x"ffffff",
   70327 => x"ffffff",
   70328 => x"ffffff",
   70329 => x"ffffff",
   70330 => x"ffffff",
   70331 => x"ffffff",
   70332 => x"ffffff",
   70333 => x"ffffff",
   70334 => x"ffffff",
   70335 => x"ffffff",
   70336 => x"ffffff",
   70337 => x"ffffff",
   70338 => x"ffffff",
   70339 => x"ffffff",
   70340 => x"ffffff",
   70341 => x"ffffff",
   70342 => x"ffffff",
   70343 => x"ffffff",
   70344 => x"ffffff",
   70345 => x"ffffff",
   70346 => x"ffffff",
   70347 => x"ffffff",
   70348 => x"ffffff",
   70349 => x"ffffff",
   70350 => x"ffffff",
   70351 => x"ffffff",
   70352 => x"ffffff",
   70353 => x"ffffff",
   70354 => x"ffffff",
   70355 => x"ffffff",
   70356 => x"ffffff",
   70357 => x"ffffff",
   70358 => x"ffffff",
   70359 => x"ffffff",
   70360 => x"ffffff",
   70361 => x"ffffff",
   70362 => x"ffffff",
   70363 => x"ffffff",
   70364 => x"ffffff",
   70365 => x"ffffff",
   70366 => x"ffffff",
   70367 => x"ffffff",
   70368 => x"ffffff",
   70369 => x"ffffff",
   70370 => x"ffffff",
   70371 => x"ffffff",
   70372 => x"ffffff",
   70373 => x"ffffff",
   70374 => x"ffffff",
   70375 => x"ffffff",
   70376 => x"ffffff",
   70377 => x"ffffff",
   70378 => x"ffffff",
   70379 => x"ffffff",
   70380 => x"ffffff",
   70381 => x"ffffff",
   70382 => x"ffffff",
   70383 => x"ffffff",
   70384 => x"ffffff",
   70385 => x"ffffff",
   70386 => x"ffffff",
   70387 => x"ffffff",
   70388 => x"ffffff",
   70389 => x"ffffff",
   70390 => x"ffffff",
   70391 => x"ffffff",
   70392 => x"ffffff",
   70393 => x"ffffff",
   70394 => x"ffffff",
   70395 => x"ffffff",
   70396 => x"ffffff",
   70397 => x"ffffff",
   70398 => x"ffffff",
   70399 => x"ffffff",
   70400 => x"ffffff",
   70401 => x"ffffff",
   70402 => x"ffffff",
   70403 => x"ffffff",
   70404 => x"ffffff",
   70405 => x"ffffff",
   70406 => x"ffffff",
   70407 => x"ffffff",
   70408 => x"ffffff",
   70409 => x"ffffff",
   70410 => x"ffffff",
   70411 => x"ffffff",
   70412 => x"ffffff",
   70413 => x"ffffff",
   70414 => x"ffffff",
   70415 => x"ffffff",
   70416 => x"ffffff",
   70417 => x"ffffff",
   70418 => x"ffffff",
   70419 => x"ffffff",
   70420 => x"ffffff",
   70421 => x"ffffff",
   70422 => x"ffffff",
   70423 => x"ffffff",
   70424 => x"ffffff",
   70425 => x"ffffff",
   70426 => x"ffffff",
   70427 => x"ffffff",
   70428 => x"ffffff",
   70429 => x"ffffff",
   70430 => x"ffffff",
   70431 => x"ffffff",
   70432 => x"ffffff",
   70433 => x"ffffff",
   70434 => x"ffffff",
   70435 => x"ffffff",
   70436 => x"ffffff",
   70437 => x"ffffff",
   70438 => x"ffffff",
   70439 => x"ffffff",
   70440 => x"ffffff",
   70441 => x"ffffff",
   70442 => x"ffffff",
   70443 => x"ffffff",
   70444 => x"ffffff",
   70445 => x"ffffff",
   70446 => x"ffffff",
   70447 => x"ffffff",
   70448 => x"ffffff",
   70449 => x"ffffff",
   70450 => x"ffffff",
   70451 => x"ffffff",
   70452 => x"ffffff",
   70453 => x"ffffff",
   70454 => x"ffffff",
   70455 => x"ffffff",
   70456 => x"ffffff",
   70457 => x"ffffff",
   70458 => x"ffffff",
   70459 => x"ffffff",
   70460 => x"ffffff",
   70461 => x"ffffff",
   70462 => x"ffffff",
   70463 => x"ffffff",
   70464 => x"ffffff",
   70465 => x"ffffff",
   70466 => x"ffffff",
   70467 => x"ffffff",
   70468 => x"ffffff",
   70469 => x"ffffff",
   70470 => x"ffffff",
   70471 => x"ffffff",
   70472 => x"ffffff",
   70473 => x"ffffff",
   70474 => x"ffffff",
   70475 => x"ffffff",
   70476 => x"ffffff",
   70477 => x"ffffff",
   70478 => x"ffffff",
   70479 => x"ffffff",
   70480 => x"ffffff",
   70481 => x"ffffff",
   70482 => x"ffffff",
   70483 => x"ffffff",
   70484 => x"ffffff",
   70485 => x"ffffff",
   70486 => x"ffffff",
   70487 => x"ffffff",
   70488 => x"ffffff",
   70489 => x"ffffff",
   70490 => x"ffffff",
   70491 => x"ffffff",
   70492 => x"ffffff",
   70493 => x"ffffff",
   70494 => x"ffffff",
   70495 => x"ffffff",
   70496 => x"ffffff",
   70497 => x"ffffff",
   70498 => x"ffffff",
   70499 => x"ffffff",
   70500 => x"ffffff",
   70501 => x"ffffff",
   70502 => x"ffffff",
   70503 => x"ffffff",
   70504 => x"ffffff",
   70505 => x"ffffff",
   70506 => x"ffffff",
   70507 => x"ffffff",
   70508 => x"ffffff",
   70509 => x"ffffff",
   70510 => x"ffffff",
   70511 => x"ffffff",
   70512 => x"ffffff",
   70513 => x"ffffff",
   70514 => x"ffffff",
   70515 => x"ffffff",
   70516 => x"ffffff",
   70517 => x"ffffff",
   70518 => x"ffffff",
   70519 => x"ffffff",
   70520 => x"ffffff",
   70521 => x"ffffff",
   70522 => x"ffffff",
   70523 => x"ffffff",
   70524 => x"ffffff",
   70525 => x"ffffff",
   70526 => x"ffffff",
   70527 => x"ffffff",
   70528 => x"ffffff",
   70529 => x"ffffff",
   70530 => x"ffffff",
   70531 => x"ffffff",
   70532 => x"ffffff",
   70533 => x"ffffff",
   70534 => x"ffffff",
   70535 => x"ffffff",
   70536 => x"ffffff",
   70537 => x"ffffff",
   70538 => x"ffffff",
   70539 => x"ffffff",
   70540 => x"ffffff",
   70541 => x"ffffff",
   70542 => x"ffffff",
   70543 => x"ffffff",
   70544 => x"ffffff",
   70545 => x"ffffff",
   70546 => x"ffffff",
   70547 => x"ffffff",
   70548 => x"ffffff",
   70549 => x"ffffff",
   70550 => x"ffffff",
   70551 => x"ffffff",
   70552 => x"ffffff",
   70553 => x"ffffff",
   70554 => x"ffffff",
   70555 => x"ffffff",
   70556 => x"ffffff",
   70557 => x"ffffff",
   70558 => x"ffffff",
   70559 => x"ffffff",
   70560 => x"ffffff",
   70561 => x"ffffff",
   70562 => x"ffffff",
   70563 => x"ffffff",
   70564 => x"ffffff",
   70565 => x"ffffff",
   70566 => x"ffffff",
   70567 => x"ffffff",
   70568 => x"ffffff",
   70569 => x"ffffff",
   70570 => x"ffffff",
   70571 => x"ffffff",
   70572 => x"ffffff",
   70573 => x"ffffff",
   70574 => x"ffffff",
   70575 => x"ffffff",
   70576 => x"ffffff",
   70577 => x"ffffff",
   70578 => x"ffffff",
   70579 => x"ffffff",
   70580 => x"ffffff",
   70581 => x"ffffff",
   70582 => x"ffffff",
   70583 => x"ffffff",
   70584 => x"ffffff",
   70585 => x"ffffff",
   70586 => x"ffffff",
   70587 => x"ffffff",
   70588 => x"ffffff",
   70589 => x"ffffff",
   70590 => x"ffffff",
   70591 => x"ffffff",
   70592 => x"ffffff",
   70593 => x"ffffff",
   70594 => x"ffffff",
   70595 => x"ffffff",
   70596 => x"ffffff",
   70597 => x"ffffff",
   70598 => x"ffffff",
   70599 => x"ffffff",
   70600 => x"ffffff",
   70601 => x"ffffff",
   70602 => x"ffffff",
   70603 => x"ffffff",
   70604 => x"ffffff",
   70605 => x"ffffff",
   70606 => x"ffffff",
   70607 => x"ffffff",
   70608 => x"ffffff",
   70609 => x"ffffff",
   70610 => x"ffffff",
   70611 => x"ffffff",
   70612 => x"ffffff",
   70613 => x"ffffff",
   70614 => x"ffffff",
   70615 => x"ffffff",
   70616 => x"ffffff",
   70617 => x"ffffff",
   70618 => x"ffffff",
   70619 => x"ffffff",
   70620 => x"ffffff",
   70621 => x"ffffff",
   70622 => x"ffffff",
   70623 => x"ffffff",
   70624 => x"ffffff",
   70625 => x"ffffff",
   70626 => x"ffffff",
   70627 => x"ffffff",
   70628 => x"ffffff",
   70629 => x"ffffff",
   70630 => x"ffffff",
   70631 => x"ffffff",
   70632 => x"ffffff",
   70633 => x"ffffff",
   70634 => x"ffffff",
   70635 => x"ffffff",
   70636 => x"ffffff",
   70637 => x"ffffff",
   70638 => x"ffffff",
   70639 => x"ffffff",
   70640 => x"ffffff",
   70641 => x"ffffff",
   70642 => x"ffffff",
   70643 => x"ffffff",
   70644 => x"ffffff",
   70645 => x"ffffff",
   70646 => x"ffffff",
   70647 => x"ffffff",
   70648 => x"ffffff",
   70649 => x"ffffff",
   70650 => x"ffffff",
   70651 => x"ffffff",
   70652 => x"ffffff",
   70653 => x"ffffff",
   70654 => x"ffffff",
   70655 => x"ffffff",
   70656 => x"ffffff",
   70657 => x"ffffff",
   70658 => x"ffffff",
   70659 => x"ffffff",
   70660 => x"ffffff",
   70661 => x"ffffff",
   70662 => x"ffffff",
   70663 => x"ffffff",
   70664 => x"ffffff",
   70665 => x"ffffff",
   70666 => x"ffffff",
   70667 => x"ffffff",
   70668 => x"ffffff",
   70669 => x"ffffff",
   70670 => x"ffffff",
   70671 => x"ffffff",
   70672 => x"ffffff",
   70673 => x"ffffff",
   70674 => x"ffffff",
   70675 => x"ffffff",
   70676 => x"ffffff",
   70677 => x"ffffff",
   70678 => x"ffffff",
   70679 => x"ffffff",
   70680 => x"ffffff",
   70681 => x"ffffff",
   70682 => x"ffffff",
   70683 => x"ffffff",
   70684 => x"ffffff",
   70685 => x"ffffff",
   70686 => x"ffffff",
   70687 => x"ffffff",
   70688 => x"ffffff",
   70689 => x"ffffff",
   70690 => x"ffffff",
   70691 => x"ffffff",
   70692 => x"ffffff",
   70693 => x"ffffff",
   70694 => x"ffffff",
   70695 => x"ffffff",
   70696 => x"ffffff",
   70697 => x"ffffff",
   70698 => x"ffffff",
   70699 => x"ffffff",
   70700 => x"ffffff",
   70701 => x"ffffff",
   70702 => x"ffffff",
   70703 => x"ffffff",
   70704 => x"ffffff",
   70705 => x"ffffff",
   70706 => x"ffffff",
   70707 => x"ffffff",
   70708 => x"ffffff",
   70709 => x"ffffff",
   70710 => x"ffffff",
   70711 => x"ffffff",
   70712 => x"ffffff",
   70713 => x"ffffff",
   70714 => x"ffffff",
   70715 => x"ffffff",
   70716 => x"ffffff",
   70717 => x"ffffff",
   70718 => x"ffffff",
   70719 => x"ffffff",
   70720 => x"ffffff",
   70721 => x"ffffff",
   70722 => x"ffffff",
   70723 => x"ffffff",
   70724 => x"ffffff",
   70725 => x"ffffff",
   70726 => x"ffffff",
   70727 => x"ffffff",
   70728 => x"ffffff",
   70729 => x"ffffff",
   70730 => x"ffffff",
   70731 => x"ffffff",
   70732 => x"ffffff",
   70733 => x"ffffff",
   70734 => x"ffffff",
   70735 => x"ffffff",
   70736 => x"ffffff",
   70737 => x"ffffff",
   70738 => x"ffffff",
   70739 => x"ffffff",
   70740 => x"ffffff",
   70741 => x"ffffff",
   70742 => x"ffffff",
   70743 => x"ffffff",
   70744 => x"ffffff",
   70745 => x"ffffff",
   70746 => x"ffffff",
   70747 => x"ffffff",
   70748 => x"ffffff",
   70749 => x"ffffff",
   70750 => x"ffffff",
   70751 => x"ffffff",
   70752 => x"ffffff",
   70753 => x"ffffff",
   70754 => x"ffffff",
   70755 => x"ffffff",
   70756 => x"ffffff",
   70757 => x"ffffff",
   70758 => x"ffffff",
   70759 => x"ffffff",
   70760 => x"ffffff",
   70761 => x"ffffff",
   70762 => x"ffffff",
   70763 => x"ffffff",
   70764 => x"ffffff",
   70765 => x"ffffff",
   70766 => x"ffffff",
   70767 => x"ffffff",
   70768 => x"ffffff",
   70769 => x"ffffff",
   70770 => x"ffffff",
   70771 => x"ffffff",
   70772 => x"ffffff",
   70773 => x"ffffff",
   70774 => x"ffffff",
   70775 => x"ffffff",
   70776 => x"ffffff",
   70777 => x"ffffff",
   70778 => x"ffffff",
   70779 => x"ffffff",
   70780 => x"ffffff",
   70781 => x"ffffff",
   70782 => x"ffffff",
   70783 => x"ffffff",
   70784 => x"ffffff",
   70785 => x"ffffff",
   70786 => x"ffffff",
   70787 => x"ffffff",
   70788 => x"ffffff",
   70789 => x"ffffff",
   70790 => x"ffffff",
   70791 => x"ffffff",
   70792 => x"ffffff",
   70793 => x"ffffff",
   70794 => x"ffffff",
   70795 => x"ffffff",
   70796 => x"ffffff",
   70797 => x"ffffff",
   70798 => x"ffffff",
   70799 => x"ffffff",
   70800 => x"ffffff",
   70801 => x"ffffff",
   70802 => x"ffffff",
   70803 => x"ffffff",
   70804 => x"ffffff",
   70805 => x"ffffff",
   70806 => x"ffffff",
   70807 => x"ffffff",
   70808 => x"ffffff",
   70809 => x"ffffff",
   70810 => x"ffffff",
   70811 => x"ffffff",
   70812 => x"ffffff",
   70813 => x"ffffff",
   70814 => x"ffffff",
   70815 => x"ffffff",
   70816 => x"ffffff",
   70817 => x"ffffff",
   70818 => x"ffffff",
   70819 => x"ffffff",
   70820 => x"ffffff",
   70821 => x"ffffff",
   70822 => x"ffffff",
   70823 => x"ffffff",
   70824 => x"ffffff",
   70825 => x"ffffff",
   70826 => x"ffffff",
   70827 => x"ffffff",
   70828 => x"ffffff",
   70829 => x"ffffff",
   70830 => x"ffffff",
   70831 => x"ffffff",
   70832 => x"ffffff",
   70833 => x"ffffff",
   70834 => x"ffffff",
   70835 => x"ffffff",
   70836 => x"ffffff",
   70837 => x"ffffff",
   70838 => x"ffffff",
   70839 => x"ffffff",
   70840 => x"ffffff",
   70841 => x"ffffff",
   70842 => x"ffffff",
   70843 => x"ffffff",
   70844 => x"ffffff",
   70845 => x"ffffff",
   70846 => x"ffffff",
   70847 => x"ffffff",
   70848 => x"ffffff",
   70849 => x"ffffff",
   70850 => x"ffffff",
   70851 => x"ffffff",
   70852 => x"ffffff",
   70853 => x"ffffff",
   70854 => x"ffffff",
   70855 => x"ffffff",
   70856 => x"ffffff",
   70857 => x"ffffff",
   70858 => x"ffffff",
   70859 => x"ffffff",
   70860 => x"ffffff",
   70861 => x"ffffff",
   70862 => x"ffffff",
   70863 => x"ffffff",
   70864 => x"ffffff",
   70865 => x"ffffff",
   70866 => x"ffffff",
   70867 => x"ffffff",
   70868 => x"ffffff",
   70869 => x"ffffff",
   70870 => x"ffffff",
   70871 => x"ffffff",
   70872 => x"ffffff",
   70873 => x"ffffff",
   70874 => x"ffffff",
   70875 => x"ffffff",
   70876 => x"ffffff",
   70877 => x"ffffff",
   70878 => x"ffffff",
   70879 => x"ffffff",
   70880 => x"ffffff",
   70881 => x"ffffff",
   70882 => x"ffffff",
   70883 => x"ffffff",
   70884 => x"ffffff",
   70885 => x"ffffff",
   70886 => x"ffffff",
   70887 => x"ffffff",
   70888 => x"ffffff",
   70889 => x"ffffff",
   70890 => x"ffffff",
   70891 => x"ffffff",
   70892 => x"ffffff",
   70893 => x"ffffff",
   70894 => x"ffffff",
   70895 => x"ffffff",
   70896 => x"ffffff",
   70897 => x"ffffff",
   70898 => x"ffffff",
   70899 => x"ffffff",
   70900 => x"ffffff",
   70901 => x"ffffff",
   70902 => x"ffffff",
   70903 => x"ffffff",
   70904 => x"ffffff",
   70905 => x"ffffff",
   70906 => x"ffffff",
   70907 => x"ffffff",
   70908 => x"ffffff",
   70909 => x"ffffff",
   70910 => x"ffffff",
   70911 => x"ffffff",
   70912 => x"ffffff",
   70913 => x"ffffff",
   70914 => x"ffffff",
   70915 => x"ffffff",
   70916 => x"ffffff",
   70917 => x"ffffff",
   70918 => x"ffffff",
   70919 => x"ffffff",
   70920 => x"ffffff",
   70921 => x"ffffff",
   70922 => x"ffffff",
   70923 => x"ffffff",
   70924 => x"ffffff",
   70925 => x"ffffff",
   70926 => x"ffffff",
   70927 => x"ffffff",
   70928 => x"ffffff",
   70929 => x"ffffff",
   70930 => x"ffffff",
   70931 => x"ffffff",
   70932 => x"ffffff",
   70933 => x"ffffff",
   70934 => x"ffffff",
   70935 => x"ffffff",
   70936 => x"ffffff",
   70937 => x"ffffff",
   70938 => x"ffffff",
   70939 => x"ffffff",
   70940 => x"ffffff",
   70941 => x"ffffff",
   70942 => x"ffffff",
   70943 => x"ffffff",
   70944 => x"ffffff",
   70945 => x"ffffff",
   70946 => x"ffffff",
   70947 => x"ffffff",
   70948 => x"ffffff",
   70949 => x"ffffff",
   70950 => x"ffffff",
   70951 => x"ffffff",
   70952 => x"ffffff",
   70953 => x"ffffff",
   70954 => x"ffffff",
   70955 => x"ffffff",
   70956 => x"ffffff",
   70957 => x"ffffff",
   70958 => x"ffffff",
   70959 => x"ffffff",
   70960 => x"ffffff",
   70961 => x"ffffff",
   70962 => x"ffffff",
   70963 => x"ffffff",
   70964 => x"ffffff",
   70965 => x"ffffff",
   70966 => x"ffffff",
   70967 => x"ffffff",
   70968 => x"ffffff",
   70969 => x"ffffff",
   70970 => x"ffffff",
   70971 => x"ffffff",
   70972 => x"ffffff",
   70973 => x"ffffff",
   70974 => x"ffffff",
   70975 => x"ffffff",
   70976 => x"ffffff",
   70977 => x"ffffff",
   70978 => x"ffffff",
   70979 => x"ffffff",
   70980 => x"ffffff",
   70981 => x"ffffff",
   70982 => x"ffffff",
   70983 => x"ffffff",
   70984 => x"ffffff",
   70985 => x"ffffff",
   70986 => x"ffffff",
   70987 => x"ffffff",
   70988 => x"ffffff",
   70989 => x"ffffff",
   70990 => x"ffffff",
   70991 => x"ffffff",
   70992 => x"ffffff",
   70993 => x"ffffff",
   70994 => x"ffffff",
   70995 => x"ffffff",
   70996 => x"ffffff",
   70997 => x"ffffff",
   70998 => x"ffffff",
   70999 => x"ffffff",
   71000 => x"ffffff",
   71001 => x"ffffff",
   71002 => x"ffffff",
   71003 => x"ffffff",
   71004 => x"ffffff",
   71005 => x"ffffff",
   71006 => x"ffffff",
   71007 => x"ffffff",
   71008 => x"ffffff",
   71009 => x"ffffff",
   71010 => x"ffffff",
   71011 => x"ffffff",
   71012 => x"ffffff",
   71013 => x"ffffff",
   71014 => x"ffffff",
   71015 => x"ffffff",
   71016 => x"ffffff",
   71017 => x"ffffff",
   71018 => x"ffffff",
   71019 => x"ffffff",
   71020 => x"ffffff",
   71021 => x"ffffff",
   71022 => x"ffffff",
   71023 => x"ffffff",
   71024 => x"ffffff",
   71025 => x"ffffff",
   71026 => x"ffffff",
   71027 => x"ffffff",
   71028 => x"ffffff",
   71029 => x"ffffff",
   71030 => x"ffffff",
   71031 => x"ffffff",
   71032 => x"ffffff",
   71033 => x"ffffff",
   71034 => x"ffffff",
   71035 => x"ffffff",
   71036 => x"ffffff",
   71037 => x"ffffff",
   71038 => x"ffffff",
   71039 => x"ffffff",
   71040 => x"ffffff",
   71041 => x"ffffff",
   71042 => x"ffffff",
   71043 => x"ffffff",
   71044 => x"ffffff",
   71045 => x"ffffff",
   71046 => x"ffffff",
   71047 => x"ffffff",
   71048 => x"ffffff",
   71049 => x"ffffff",
   71050 => x"ffffff",
   71051 => x"ffffff",
   71052 => x"ffffff",
   71053 => x"ffffff",
   71054 => x"ffffff",
   71055 => x"ffffff",
   71056 => x"ffffff",
   71057 => x"ffffff",
   71058 => x"ffffff",
   71059 => x"ffffff",
   71060 => x"ffffff",
   71061 => x"ffffff",
   71062 => x"ffffff",
   71063 => x"ffffff",
   71064 => x"ffffff",
   71065 => x"ffffff",
   71066 => x"ffffff",
   71067 => x"ffffff",
   71068 => x"ffffff",
   71069 => x"ffffff",
   71070 => x"ffffff",
   71071 => x"ffffff",
   71072 => x"ffffff",
   71073 => x"ffffff",
   71074 => x"ffffff",
   71075 => x"ffffff",
   71076 => x"ffffff",
   71077 => x"ffffff",
   71078 => x"ffffff",
   71079 => x"ffffff",
   71080 => x"ffffff",
   71081 => x"ffffff",
   71082 => x"ffffff",
   71083 => x"ffffff",
   71084 => x"ffffff",
   71085 => x"ffffff",
   71086 => x"ffffff",
   71087 => x"ffffff",
   71088 => x"ffffff",
   71089 => x"ffffff",
   71090 => x"ffffff",
   71091 => x"ffffff",
   71092 => x"ffffff",
   71093 => x"ffffff",
   71094 => x"ffffff",
   71095 => x"ffffff",
   71096 => x"ffffff",
   71097 => x"ffffff",
   71098 => x"ffffff",
   71099 => x"ffffff",
   71100 => x"ffffff",
   71101 => x"ffffff",
   71102 => x"ffffff",
   71103 => x"ffffff",
   71104 => x"ffffff",
   71105 => x"ffffff",
   71106 => x"ffffff",
   71107 => x"ffffff",
   71108 => x"ffffff",
   71109 => x"ffffff",
   71110 => x"ffffff",
   71111 => x"ffffff",
   71112 => x"ffffff",
   71113 => x"ffffff",
   71114 => x"ffffff",
   71115 => x"ffffff",
   71116 => x"ffffff",
   71117 => x"ffffff",
   71118 => x"ffffff",
   71119 => x"ffffff",
   71120 => x"ffffff",
   71121 => x"ffffff",
   71122 => x"ffffff",
   71123 => x"ffffff",
   71124 => x"ffffff",
   71125 => x"ffffff",
   71126 => x"ffffff",
   71127 => x"ffffff",
   71128 => x"ffffff",
   71129 => x"ffffff",
   71130 => x"ffffff",
   71131 => x"ffffff",
   71132 => x"ffffff",
   71133 => x"ffffff",
   71134 => x"ffffff",
   71135 => x"ffffff",
   71136 => x"ffffff",
   71137 => x"ffffff",
   71138 => x"ffffff",
   71139 => x"ffffff",
   71140 => x"ffffff",
   71141 => x"ffffff",
   71142 => x"ffffff",
   71143 => x"ffffff",
   71144 => x"ffffff",
   71145 => x"ffffff",
   71146 => x"ffffff",
   71147 => x"ffffff",
   71148 => x"ffffff",
   71149 => x"ffffff",
   71150 => x"ffffff",
   71151 => x"ffffff",
   71152 => x"ffffff",
   71153 => x"ffffff",
   71154 => x"ffffff",
   71155 => x"ffffff",
   71156 => x"ffffff",
   71157 => x"ffffff",
   71158 => x"ffffff",
   71159 => x"ffffff",
   71160 => x"ffffff",
   71161 => x"ffffff",
   71162 => x"ffffff",
   71163 => x"ffffff",
   71164 => x"ffffff",
   71165 => x"ffffff",
   71166 => x"ffffff",
   71167 => x"ffffff",
   71168 => x"ffffff",
   71169 => x"ffffff",
   71170 => x"ffffff",
   71171 => x"ffffff",
   71172 => x"ffffff",
   71173 => x"ffffff",
   71174 => x"ffffff",
   71175 => x"ffffff",
   71176 => x"ffffff",
   71177 => x"ffffff",
   71178 => x"ffffff",
   71179 => x"ffffff",
   71180 => x"ffffff",
   71181 => x"ffffff",
   71182 => x"ffffff",
   71183 => x"ffffff",
   71184 => x"ffffff",
   71185 => x"ffffff",
   71186 => x"ffffff",
   71187 => x"ffffff",
   71188 => x"ffffff",
   71189 => x"ffffff",
   71190 => x"ffffff",
   71191 => x"ffffff",
   71192 => x"ffffff",
   71193 => x"ffffff",
   71194 => x"ffffff",
   71195 => x"ffffff",
   71196 => x"ffffff",
   71197 => x"ffffff",
   71198 => x"ffffff",
   71199 => x"ffffff",
   71200 => x"ffffff",
   71201 => x"ffffff",
   71202 => x"ffffff",
   71203 => x"ffffff",
   71204 => x"ffffff",
   71205 => x"ffffff",
   71206 => x"ffffff",
   71207 => x"ffffff",
   71208 => x"ffffff",
   71209 => x"ffffff",
   71210 => x"ffffff",
   71211 => x"ffffff",
   71212 => x"ffffff",
   71213 => x"ffffff",
   71214 => x"ffffff",
   71215 => x"ffffff",
   71216 => x"ffffff",
   71217 => x"ffffff",
   71218 => x"ffffff",
   71219 => x"ffffff",
   71220 => x"ffffff",
   71221 => x"ffffff",
   71222 => x"ffffff",
   71223 => x"ffffff",
   71224 => x"ffffff",
   71225 => x"ffffff",
   71226 => x"ffffff",
   71227 => x"ffffff",
   71228 => x"ffffff",
   71229 => x"ffffff",
   71230 => x"ffffff",
   71231 => x"ffffff",
   71232 => x"ffffff",
   71233 => x"ffffff",
   71234 => x"ffffff",
   71235 => x"ffffff",
   71236 => x"ffffff",
   71237 => x"ffffff",
   71238 => x"ffffff",
   71239 => x"ffffff",
   71240 => x"ffffff",
   71241 => x"ffffff",
   71242 => x"ffffff",
   71243 => x"ffffff",
   71244 => x"ffffff",
   71245 => x"ffffff",
   71246 => x"ffffff",
   71247 => x"ffffff",
   71248 => x"ffffff",
   71249 => x"ffffff",
   71250 => x"ffffff",
   71251 => x"ffffff",
   71252 => x"ffffff",
   71253 => x"ffffff",
   71254 => x"ffffff",
   71255 => x"ffffff",
   71256 => x"ffffff",
   71257 => x"ffffff",
   71258 => x"ffffff",
   71259 => x"ffffff",
   71260 => x"ffffff",
   71261 => x"ffffff",
   71262 => x"ffffff",
   71263 => x"ffffff",
   71264 => x"ffffff",
   71265 => x"ffffff",
   71266 => x"ffffff",
   71267 => x"ffffff",
   71268 => x"ffffff",
   71269 => x"ffffff",
   71270 => x"ffffff",
   71271 => x"ffffff",
   71272 => x"ffffff",
   71273 => x"ffffff",
   71274 => x"ffffff",
   71275 => x"ffffff",
   71276 => x"ffffff",
   71277 => x"ffffff",
   71278 => x"ffffff",
   71279 => x"ffffff",
   71280 => x"ffffff",
   71281 => x"ffffff",
   71282 => x"ffffff",
   71283 => x"ffffff",
   71284 => x"ffffff",
   71285 => x"ffffff",
   71286 => x"ffffff",
   71287 => x"ffffff",
   71288 => x"ffffff",
   71289 => x"ffffff",
   71290 => x"ffffff",
   71291 => x"ffffff",
   71292 => x"ffffff",
   71293 => x"ffffff",
   71294 => x"ffffff",
   71295 => x"ffffff",
   71296 => x"ffffff",
   71297 => x"ffffff",
   71298 => x"ffffff",
   71299 => x"ffffff",
   71300 => x"ffffff",
   71301 => x"ffffff",
   71302 => x"ffffff",
   71303 => x"ffffff",
   71304 => x"ffffff",
   71305 => x"ffffff",
   71306 => x"ffffff",
   71307 => x"ffffff",
   71308 => x"ffffff",
   71309 => x"ffffff",
   71310 => x"ffffff",
   71311 => x"ffffff",
   71312 => x"ffffff",
   71313 => x"ffffff",
   71314 => x"ffffff",
   71315 => x"ffffff",
   71316 => x"ffffff",
   71317 => x"ffffff",
   71318 => x"ffffff",
   71319 => x"ffffff",
   71320 => x"ffffff",
   71321 => x"ffffff",
   71322 => x"ffffff",
   71323 => x"ffffff",
   71324 => x"ffffff",
   71325 => x"ffffff",
   71326 => x"ffffff",
   71327 => x"ffffff",
   71328 => x"ffffff",
   71329 => x"ffffff",
   71330 => x"ffffff",
   71331 => x"ffffff",
   71332 => x"ffffff",
   71333 => x"ffffff",
   71334 => x"ffffff",
   71335 => x"ffffff",
   71336 => x"ffffff",
   71337 => x"ffffff",
   71338 => x"ffffff",
   71339 => x"ffffff",
   71340 => x"ffffff",
   71341 => x"ffffff",
   71342 => x"ffffff",
   71343 => x"ffffff",
   71344 => x"ffffff",
   71345 => x"ffffff",
   71346 => x"ffffff",
   71347 => x"ffffff",
   71348 => x"ffffff",
   71349 => x"ffffff",
   71350 => x"ffffff",
   71351 => x"ffffff",
   71352 => x"ffffff",
   71353 => x"ffffff",
   71354 => x"ffffff",
   71355 => x"ffffff",
   71356 => x"ffffff",
   71357 => x"ffffff",
   71358 => x"ffffff",
   71359 => x"ffffff",
   71360 => x"ffffff",
   71361 => x"ffffff",
   71362 => x"ffffff",
   71363 => x"ffffff",
   71364 => x"ffffff",
   71365 => x"ffffff",
   71366 => x"ffffff",
   71367 => x"ffffff",
   71368 => x"ffffff",
   71369 => x"ffffff",
   71370 => x"ffffff",
   71371 => x"ffffff",
   71372 => x"ffffff",
   71373 => x"ffffff",
   71374 => x"ffffff",
   71375 => x"ffffff",
   71376 => x"ffffff",
   71377 => x"ffffff",
   71378 => x"ffffff",
   71379 => x"ffffff",
   71380 => x"ffffff",
   71381 => x"ffffff",
   71382 => x"ffffff",
   71383 => x"ffffff",
   71384 => x"ffffff",
   71385 => x"ffffff",
   71386 => x"ffffff",
   71387 => x"ffffff",
   71388 => x"ffffff",
   71389 => x"ffffff",
   71390 => x"ffffff",
   71391 => x"ffffff",
   71392 => x"ffffff",
   71393 => x"ffffff",
   71394 => x"ffffff",
   71395 => x"ffffff",
   71396 => x"ffffff",
   71397 => x"ffffff",
   71398 => x"ffffff",
   71399 => x"ffffff",
   71400 => x"ffffff",
   71401 => x"ffffff",
   71402 => x"ffffff",
   71403 => x"ffffff",
   71404 => x"ffffff",
   71405 => x"ffffff",
   71406 => x"ffffff",
   71407 => x"ffffff",
   71408 => x"ffffff",
   71409 => x"ffffff",
   71410 => x"ffffff",
   71411 => x"ffffff",
   71412 => x"ffffff",
   71413 => x"ffffff",
   71414 => x"ffffff",
   71415 => x"ffffff",
   71416 => x"ffffff",
   71417 => x"ffffff",
   71418 => x"ffffff",
   71419 => x"ffffff",
   71420 => x"ffffff",
   71421 => x"ffffff",
   71422 => x"ffffff",
   71423 => x"ffffff",
   71424 => x"ffffff",
   71425 => x"ffffff",
   71426 => x"ffffff",
   71427 => x"ffffff",
   71428 => x"ffffff",
   71429 => x"ffffff",
   71430 => x"ffffff",
   71431 => x"ffffff",
   71432 => x"ffffff",
   71433 => x"ffffff",
   71434 => x"ffffff",
   71435 => x"ffffff",
   71436 => x"ffffff",
   71437 => x"ffffff",
   71438 => x"ffffff",
   71439 => x"ffffff",
   71440 => x"ffffff",
   71441 => x"ffffff",
   71442 => x"ffffff",
   71443 => x"ffffff",
   71444 => x"ffffff",
   71445 => x"ffffff",
   71446 => x"ffffff",
   71447 => x"ffffff",
   71448 => x"ffffff",
   71449 => x"ffffff",
   71450 => x"ffffff",
   71451 => x"ffffff",
   71452 => x"ffffff",
   71453 => x"ffffff",
   71454 => x"ffffff",
   71455 => x"ffffff",
   71456 => x"ffffff",
   71457 => x"ffffff",
   71458 => x"ffffff",
   71459 => x"ffffff",
   71460 => x"ffffff",
   71461 => x"ffffff",
   71462 => x"ffffff",
   71463 => x"ffffff",
   71464 => x"ffffff",
   71465 => x"ffffff",
   71466 => x"ffffff",
   71467 => x"ffffff",
   71468 => x"ffffff",
   71469 => x"ffffff",
   71470 => x"ffffff",
   71471 => x"ffffff",
   71472 => x"ffffff",
   71473 => x"ffffff",
   71474 => x"ffffff",
   71475 => x"ffffff",
   71476 => x"ffffff",
   71477 => x"ffffff",
   71478 => x"ffffff",
   71479 => x"ffffff",
   71480 => x"ffffff",
   71481 => x"ffffff",
   71482 => x"ffffff",
   71483 => x"ffffff",
   71484 => x"ffffff",
   71485 => x"ffffff",
   71486 => x"ffffff",
   71487 => x"ffffff",
   71488 => x"ffffff",
   71489 => x"ffffff",
   71490 => x"ffffff",
   71491 => x"ffffff",
   71492 => x"ffffff",
   71493 => x"ffffff",
   71494 => x"ffffff",
   71495 => x"ffffff",
   71496 => x"ffffff",
   71497 => x"ffffff",
   71498 => x"ffffff",
   71499 => x"ffffff",
   71500 => x"ffffff",
   71501 => x"ffffff",
   71502 => x"ffffff",
   71503 => x"ffffff",
   71504 => x"ffffff",
   71505 => x"ffffff",
   71506 => x"ffffff",
   71507 => x"ffffff",
   71508 => x"ffffff",
   71509 => x"ffffff",
   71510 => x"ffffff",
   71511 => x"ffffff",
   71512 => x"ffffff",
   71513 => x"ffffff",
   71514 => x"ffffff",
   71515 => x"ffffff",
   71516 => x"ffffff",
   71517 => x"ffffff",
   71518 => x"ffffff",
   71519 => x"ffffff",
   71520 => x"ffffff",
   71521 => x"ffffff",
   71522 => x"ffffff",
   71523 => x"ffffff",
   71524 => x"ffffff",
   71525 => x"ffffff",
   71526 => x"ffffff",
   71527 => x"ffffff",
   71528 => x"ffffff",
   71529 => x"ffffff",
   71530 => x"ffffff",
   71531 => x"ffffff",
   71532 => x"ffffff",
   71533 => x"ffffff",
   71534 => x"ffffff",
   71535 => x"ffffff",
   71536 => x"ffffff",
   71537 => x"ffffff",
   71538 => x"ffffff",
   71539 => x"ffffff",
   71540 => x"ffffff",
   71541 => x"ffffff",
   71542 => x"ffffff",
   71543 => x"ffffff",
   71544 => x"ffffff",
   71545 => x"ffffff",
   71546 => x"ffffff",
   71547 => x"ffffff",
   71548 => x"ffffff",
   71549 => x"ffffff",
   71550 => x"ffffff",
   71551 => x"ffffff",
   71552 => x"ffffff",
   71553 => x"ffffff",
   71554 => x"ffffff",
   71555 => x"ffffff",
   71556 => x"ffffff",
   71557 => x"ffffff",
   71558 => x"ffffff",
   71559 => x"ffffff",
   71560 => x"ffffff",
   71561 => x"ffffff",
   71562 => x"ffffff",
   71563 => x"ffffff",
   71564 => x"ffffff",
   71565 => x"ffffff",
   71566 => x"ffffff",
   71567 => x"ffffff",
   71568 => x"ffffff",
   71569 => x"ffffff",
   71570 => x"ffffff",
   71571 => x"ffffff",
   71572 => x"ffffff",
   71573 => x"ffffff",
   71574 => x"ffffff",
   71575 => x"ffffff",
   71576 => x"ffffff",
   71577 => x"ffffff",
   71578 => x"ffffff",
   71579 => x"ffffff",
   71580 => x"ffffff",
   71581 => x"ffffff",
   71582 => x"ffffff",
   71583 => x"ffffff",
   71584 => x"ffffff",
   71585 => x"ffffff",
   71586 => x"ffffff",
   71587 => x"ffffff",
   71588 => x"ffffff",
   71589 => x"ffffff",
   71590 => x"ffffff",
   71591 => x"ffffff",
   71592 => x"ffffff",
   71593 => x"ffffff",
   71594 => x"ffffff",
   71595 => x"ffffff",
   71596 => x"ffffff",
   71597 => x"ffffff",
   71598 => x"ffffff",
   71599 => x"ffffff",
   71600 => x"ffffff",
   71601 => x"ffffff",
   71602 => x"ffffff",
   71603 => x"ffffff",
   71604 => x"ffffff",
   71605 => x"ffffff",
   71606 => x"ffffff",
   71607 => x"ffffff",
   71608 => x"ffffff",
   71609 => x"ffffff",
   71610 => x"ffffff",
   71611 => x"ffffff",
   71612 => x"ffffff",
   71613 => x"ffffff",
   71614 => x"ffffff",
   71615 => x"ffffff",
   71616 => x"ffffff",
   71617 => x"ffffff",
   71618 => x"ffffff",
   71619 => x"ffffff",
   71620 => x"ffffff",
   71621 => x"ffffff",
   71622 => x"ffffff",
   71623 => x"ffffff",
   71624 => x"ffffff",
   71625 => x"ffffff",
   71626 => x"ffffff",
   71627 => x"ffffff",
   71628 => x"ffffff",
   71629 => x"ffffff",
   71630 => x"ffffff",
   71631 => x"ffffff",
   71632 => x"ffffff",
   71633 => x"ffffff",
   71634 => x"ffffff",
   71635 => x"ffffff",
   71636 => x"ffffff",
   71637 => x"ffffff",
   71638 => x"ffffff",
   71639 => x"ffffff",
   71640 => x"ffffff",
   71641 => x"ffffff",
   71642 => x"ffffff",
   71643 => x"ffffff",
   71644 => x"ffffff",
   71645 => x"ffffff",
   71646 => x"ffffff",
   71647 => x"ffffff",
   71648 => x"ffffff",
   71649 => x"ffffff",
   71650 => x"ffffff",
   71651 => x"ffffff",
   71652 => x"ffffff",
   71653 => x"ffffff",
   71654 => x"ffffff",
   71655 => x"ffffff",
   71656 => x"ffffff",
   71657 => x"ffffff",
   71658 => x"ffffff",
   71659 => x"ffffff",
   71660 => x"ffffff",
   71661 => x"ffffff",
   71662 => x"ffffff",
   71663 => x"ffffff",
   71664 => x"ffffff",
   71665 => x"ffffff",
   71666 => x"ffffff",
   71667 => x"ffffff",
   71668 => x"ffffff",
   71669 => x"ffffff",
   71670 => x"ffffff",
   71671 => x"ffffff",
   71672 => x"ffffff",
   71673 => x"ffffff",
   71674 => x"ffffff",
   71675 => x"ffffff",
   71676 => x"ffffff",
   71677 => x"ffffff",
   71678 => x"ffffff",
   71679 => x"ffffff",
   71680 => x"ffffff",
   71681 => x"ffffff",
   71682 => x"ffffff",
   71683 => x"ffffff",
   71684 => x"ffffff",
   71685 => x"ffffff",
   71686 => x"ffffff",
   71687 => x"ffffff",
   71688 => x"ffffff",
   71689 => x"ffffff",
   71690 => x"ffffff",
   71691 => x"ffffff",
   71692 => x"ffffff",
   71693 => x"ffffff",
   71694 => x"ffffff",
   71695 => x"ffffff",
   71696 => x"ffffff",
   71697 => x"ffffff",
   71698 => x"ffffff",
   71699 => x"ffffff",
   71700 => x"ffffff",
   71701 => x"ffffff",
   71702 => x"ffffff",
   71703 => x"ffffff",
   71704 => x"ffffff",
   71705 => x"ffffff",
   71706 => x"ffffff",
   71707 => x"ffffff",
   71708 => x"ffffff",
   71709 => x"ffffff",
   71710 => x"ffffff",
   71711 => x"ffffff",
   71712 => x"ffffff",
   71713 => x"ffffff",
   71714 => x"ffffff",
   71715 => x"ffffff",
   71716 => x"ffffff",
   71717 => x"ffffff",
   71718 => x"ffffff",
   71719 => x"ffffff",
   71720 => x"ffffff",
   71721 => x"ffffff",
   71722 => x"ffffff",
   71723 => x"ffffff",
   71724 => x"ffffff",
   71725 => x"ffffff",
   71726 => x"ffffff",
   71727 => x"ffffff",
   71728 => x"ffffff",
   71729 => x"ffffff",
   71730 => x"ffffff",
   71731 => x"ffffff",
   71732 => x"ffffff",
   71733 => x"ffffff",
   71734 => x"ffffff",
   71735 => x"ffffff",
   71736 => x"ffffff",
   71737 => x"ffffff",
   71738 => x"ffffff",
   71739 => x"ffffff",
   71740 => x"ffffff",
   71741 => x"ffffff",
   71742 => x"ffffff",
   71743 => x"ffffff",
   71744 => x"ffffff",
   71745 => x"ffffff",
   71746 => x"ffffff",
   71747 => x"ffffff",
   71748 => x"ffffff",
   71749 => x"ffffff",
   71750 => x"ffffff",
   71751 => x"ffffff",
   71752 => x"ffffff",
   71753 => x"ffffff",
   71754 => x"ffffff",
   71755 => x"ffffff",
   71756 => x"ffffff",
   71757 => x"ffffff",
   71758 => x"ffffff",
   71759 => x"ffffff",
   71760 => x"ffffff",
   71761 => x"ffffff",
   71762 => x"ffffff",
   71763 => x"ffffff",
   71764 => x"ffffff",
   71765 => x"ffffff",
   71766 => x"ffffff",
   71767 => x"ffffff",
   71768 => x"ffffff",
   71769 => x"ffffff",
   71770 => x"ffffff",
   71771 => x"ffffff",
   71772 => x"ffffff",
   71773 => x"ffffff",
   71774 => x"ffffff",
   71775 => x"ffffff",
   71776 => x"ffffff",
   71777 => x"ffffff",
   71778 => x"ffffff",
   71779 => x"ffffff",
   71780 => x"ffffff",
   71781 => x"ffffff",
   71782 => x"ffffff",
   71783 => x"ffffff",
   71784 => x"ffffff",
   71785 => x"ffffff",
   71786 => x"ffffff",
   71787 => x"ffffff",
   71788 => x"ffffff",
   71789 => x"ffffff",
   71790 => x"ffffff",
   71791 => x"ffffff",
   71792 => x"ffffff",
   71793 => x"ffffff",
   71794 => x"ffffff",
   71795 => x"ffffff",
   71796 => x"ffffff",
   71797 => x"ffffff",
   71798 => x"ffffff",
   71799 => x"ffffff",
   71800 => x"ffffff",
   71801 => x"ffffff",
   71802 => x"ffffff",
   71803 => x"ffffff",
   71804 => x"ffffff",
   71805 => x"ffffff",
   71806 => x"ffffff",
   71807 => x"ffffff",
   71808 => x"ffffff",
   71809 => x"ffffff",
   71810 => x"ffffff",
   71811 => x"ffffff",
   71812 => x"ffffff",
   71813 => x"ffffff",
   71814 => x"ffffff",
   71815 => x"ffffff",
   71816 => x"ffffff",
   71817 => x"ffffff",
   71818 => x"ffffff",
   71819 => x"ffffff",
   71820 => x"ffffff",
   71821 => x"ffffff",
   71822 => x"ffffff",
   71823 => x"ffffff",
   71824 => x"ffffff",
   71825 => x"ffffff",
   71826 => x"ffffff",
   71827 => x"ffffff",
   71828 => x"ffffff",
   71829 => x"ffffff",
   71830 => x"ffffff",
   71831 => x"ffffff",
   71832 => x"ffffff",
   71833 => x"ffffff",
   71834 => x"ffffff",
   71835 => x"ffffff",
   71836 => x"ffffff",
   71837 => x"ffffff",
   71838 => x"ffffff",
   71839 => x"ffffff",
   71840 => x"ffffff",
   71841 => x"ffffff",
   71842 => x"ffffff",
   71843 => x"ffffff",
   71844 => x"ffffff",
   71845 => x"ffffff",
   71846 => x"ffffff",
   71847 => x"ffffff",
   71848 => x"ffffff",
   71849 => x"ffffff",
   71850 => x"ffffff",
   71851 => x"ffffff",
   71852 => x"ffffff",
   71853 => x"ffffff",
   71854 => x"ffffff",
   71855 => x"ffffff",
   71856 => x"ffffff",
   71857 => x"ffffff",
   71858 => x"ffffff",
   71859 => x"ffffff",
   71860 => x"ffffff",
   71861 => x"ffffff",
   71862 => x"ffffff",
   71863 => x"ffffff",
   71864 => x"ffffff",
   71865 => x"ffffff",
   71866 => x"ffffff",
   71867 => x"ffffff",
   71868 => x"ffffff",
   71869 => x"ffffff",
   71870 => x"ffffff",
   71871 => x"ffffff",
   71872 => x"ffffff",
   71873 => x"ffffff",
   71874 => x"ffffff",
   71875 => x"ffffff",
   71876 => x"ffffff",
   71877 => x"ffffff",
   71878 => x"ffffff",
   71879 => x"ffffff",
   71880 => x"ffffff",
   71881 => x"ffffff",
   71882 => x"ffffff",
   71883 => x"ffffff",
   71884 => x"ffffff",
   71885 => x"ffffff",
   71886 => x"ffffff",
   71887 => x"ffffff",
   71888 => x"ffffff",
   71889 => x"ffffff",
   71890 => x"ffffff",
   71891 => x"ffffff",
   71892 => x"ffffff",
   71893 => x"ffffff",
   71894 => x"ffffff",
   71895 => x"ffffff",
   71896 => x"ffffff",
   71897 => x"ffffff",
   71898 => x"ffffff",
   71899 => x"ffffff",
   71900 => x"ffffff",
   71901 => x"ffffff",
   71902 => x"ffffff",
   71903 => x"ffffff",
   71904 => x"ffffff",
   71905 => x"ffffff",
   71906 => x"ffffff",
   71907 => x"ffffff",
   71908 => x"ffffff",
   71909 => x"ffffff",
   71910 => x"ffffff",
   71911 => x"ffffff",
   71912 => x"ffffff",
   71913 => x"ffffff",
   71914 => x"ffffff",
   71915 => x"ffffff",
   71916 => x"ffffff",
   71917 => x"ffffff",
   71918 => x"ffffff",
   71919 => x"ffffff",
   71920 => x"ffffff",
   71921 => x"ffffff",
   71922 => x"ffffff",
   71923 => x"ffffff",
   71924 => x"ffffff",
   71925 => x"ffffff",
   71926 => x"ffffff",
   71927 => x"ffffff",
   71928 => x"ffffff",
   71929 => x"ffffff",
   71930 => x"ffffff",
   71931 => x"ffffff",
   71932 => x"ffffff",
   71933 => x"ffffff",
   71934 => x"ffffff",
   71935 => x"ffffff",
   71936 => x"ffffff",
   71937 => x"ffffff",
   71938 => x"ffffff",
   71939 => x"ffffff",
   71940 => x"ffffff",
   71941 => x"ffffff",
   71942 => x"ffffff",
   71943 => x"ffffff",
   71944 => x"ffffff",
   71945 => x"ffffff",
   71946 => x"ffffff",
   71947 => x"ffffff",
   71948 => x"ffffff",
   71949 => x"ffffff",
   71950 => x"ffffff",
   71951 => x"ffffff",
   71952 => x"ffffff",
   71953 => x"ffffff",
   71954 => x"ffffff",
   71955 => x"ffffff",
   71956 => x"ffffff",
   71957 => x"ffffff",
   71958 => x"ffffff",
   71959 => x"ffffff",
   71960 => x"ffffff",
   71961 => x"ffffff",
   71962 => x"ffffff",
   71963 => x"ffffff",
   71964 => x"ffffff",
   71965 => x"ffffff",
   71966 => x"ffffff",
   71967 => x"ffffff",
   71968 => x"ffffff",
   71969 => x"ffffff",
   71970 => x"ffffff",
   71971 => x"ffffff",
   71972 => x"ffffff",
   71973 => x"ffffff",
   71974 => x"ffffff",
   71975 => x"ffffff",
   71976 => x"ffffff",
   71977 => x"ffffff",
   71978 => x"ffffff",
   71979 => x"ffffff",
   71980 => x"ffffff",
   71981 => x"ffffff",
   71982 => x"ffffff",
   71983 => x"ffffff",
   71984 => x"ffffff",
   71985 => x"ffffff",
   71986 => x"ffffff",
   71987 => x"ffffff",
   71988 => x"ffffff",
   71989 => x"ffffff",
   71990 => x"ffffff",
   71991 => x"ffffff",
   71992 => x"ffffff",
   71993 => x"ffffff",
   71994 => x"ffffff",
   71995 => x"ffffff",
   71996 => x"ffffff",
   71997 => x"ffffff",
   71998 => x"ffffff",
   71999 => x"ffffff",
   72000 => x"ffffff",
   72001 => x"ffffff",
   72002 => x"ffffff",
   72003 => x"ffffff",
   72004 => x"ffffff",
   72005 => x"ffffff",
   72006 => x"ffffff",
   72007 => x"ffffff",
   72008 => x"ffffff",
   72009 => x"ffffff",
   72010 => x"ffffff",
   72011 => x"ffffff",
   72012 => x"ffffff",
   72013 => x"ffffff",
   72014 => x"ffffff",
   72015 => x"ffffff",
   72016 => x"ffffff",
   72017 => x"ffffff",
   72018 => x"ffffff",
   72019 => x"ffffff",
   72020 => x"ffffff",
   72021 => x"ffffff",
   72022 => x"ffffff",
   72023 => x"ffffff",
   72024 => x"ffffff",
   72025 => x"ffffff",
   72026 => x"ffffff",
   72027 => x"ffffff",
   72028 => x"ffffff",
   72029 => x"ffffff",
   72030 => x"ffffff",
   72031 => x"ffffff",
   72032 => x"ffffff",
   72033 => x"ffffff",
   72034 => x"ffffff",
   72035 => x"ffffff",
   72036 => x"ffffff",
   72037 => x"ffffff",
   72038 => x"ffffff",
   72039 => x"ffffff",
   72040 => x"ffffff",
   72041 => x"ffffff",
   72042 => x"ffffff",
   72043 => x"ffffff",
   72044 => x"ffffff",
   72045 => x"ffffff",
   72046 => x"ffffff",
   72047 => x"ffffff",
   72048 => x"ffffff",
   72049 => x"ffffff",
   72050 => x"ffffff",
   72051 => x"ffffff",
   72052 => x"ffffff",
   72053 => x"ffffff",
   72054 => x"ffffff",
   72055 => x"ffffff",
   72056 => x"ffffff",
   72057 => x"ffffff",
   72058 => x"ffffff",
   72059 => x"ffffff",
   72060 => x"ffffff",
   72061 => x"ffffff",
   72062 => x"ffffff",
   72063 => x"ffffff",
   72064 => x"ffffff",
   72065 => x"ffffff",
   72066 => x"ffffff",
   72067 => x"ffffff",
   72068 => x"ffffff",
   72069 => x"ffffff",
   72070 => x"ffffff",
   72071 => x"ffffff",
   72072 => x"ffffff",
   72073 => x"ffffff",
   72074 => x"ffffff",
   72075 => x"ffffff",
   72076 => x"ffffff",
   72077 => x"ffffff",
   72078 => x"ffffff",
   72079 => x"ffffff",
   72080 => x"ffffff",
   72081 => x"ffffff",
   72082 => x"ffffff",
   72083 => x"ffffff",
   72084 => x"ffffff",
   72085 => x"ffffff",
   72086 => x"ffffff",
   72087 => x"ffffff",
   72088 => x"ffffff",
   72089 => x"ffffff",
   72090 => x"ffffff",
   72091 => x"ffffff",
   72092 => x"ffffff",
   72093 => x"ffffff",
   72094 => x"ffffff",
   72095 => x"ffffff",
   72096 => x"ffffff",
   72097 => x"ffffff",
   72098 => x"ffffff",
   72099 => x"ffffff",
   72100 => x"ffffff",
   72101 => x"ffffff",
   72102 => x"ffffff",
   72103 => x"ffffff",
   72104 => x"ffffff",
   72105 => x"ffffff",
   72106 => x"ffffff",
   72107 => x"ffffff",
   72108 => x"ffffff",
   72109 => x"ffffff",
   72110 => x"ffffff",
   72111 => x"ffffff",
   72112 => x"ffffff",
   72113 => x"ffffff",
   72114 => x"ffffff",
   72115 => x"ffffff",
   72116 => x"ffffff",
   72117 => x"ffffff",
   72118 => x"ffffff",
   72119 => x"ffffff",
   72120 => x"ffffff",
   72121 => x"ffffff",
   72122 => x"ffffff",
   72123 => x"ffffff",
   72124 => x"ffffff",
   72125 => x"ffffff",
   72126 => x"ffffff",
   72127 => x"ffffff",
   72128 => x"ffffff",
   72129 => x"ffffff",
   72130 => x"ffffff",
   72131 => x"ffffff",
   72132 => x"ffffff",
   72133 => x"ffffff",
   72134 => x"ffffff",
   72135 => x"ffffff",
   72136 => x"ffffff",
   72137 => x"ffffff",
   72138 => x"ffffff",
   72139 => x"ffffff",
   72140 => x"ffffff",
   72141 => x"ffffff",
   72142 => x"ffffff",
   72143 => x"ffffff",
   72144 => x"ffffff",
   72145 => x"ffffff",
   72146 => x"ffffff",
   72147 => x"ffffff",
   72148 => x"ffffff",
   72149 => x"ffffff",
   72150 => x"ffffff",
   72151 => x"ffffff",
   72152 => x"ffffff",
   72153 => x"ffffff",
   72154 => x"ffffff",
   72155 => x"ffffff",
   72156 => x"ffffff",
   72157 => x"ffffff",
   72158 => x"ffffff",
   72159 => x"ffffff",
   72160 => x"ffffff",
   72161 => x"ffffff",
   72162 => x"ffffff",
   72163 => x"ffffff",
   72164 => x"ffffff",
   72165 => x"ffffff",
   72166 => x"ffffff",
   72167 => x"ffffff",
   72168 => x"ffffff",
   72169 => x"ffffff",
   72170 => x"ffffff",
   72171 => x"ffffff",
   72172 => x"ffffff",
   72173 => x"ffffff",
   72174 => x"ffffff",
   72175 => x"ffffff",
   72176 => x"ffffff",
   72177 => x"ffffff",
   72178 => x"ffffff",
   72179 => x"ffffff",
   72180 => x"ffffff",
   72181 => x"ffffff",
   72182 => x"ffffff",
   72183 => x"ffffff",
   72184 => x"ffffff",
   72185 => x"ffffff",
   72186 => x"ffffff",
   72187 => x"ffffff",
   72188 => x"ffffff",
   72189 => x"ffffff",
   72190 => x"ffffff",
   72191 => x"ffffff",
   72192 => x"ffffff",
   72193 => x"ffffff",
   72194 => x"ffffff",
   72195 => x"ffffff",
   72196 => x"ffffff",
   72197 => x"ffffff",
   72198 => x"ffffff",
   72199 => x"ffffff",
   72200 => x"ffffff",
   72201 => x"ffffff",
   72202 => x"ffffff",
   72203 => x"ffffff",
   72204 => x"ffffff",
   72205 => x"ffffff",
   72206 => x"ffffff",
   72207 => x"ffffff",
   72208 => x"ffffff",
   72209 => x"ffffff",
   72210 => x"ffffff",
   72211 => x"ffffff",
   72212 => x"ffffff",
   72213 => x"ffffff",
   72214 => x"ffffff",
   72215 => x"ffffff",
   72216 => x"ffffff",
   72217 => x"ffffff",
   72218 => x"ffffff",
   72219 => x"ffffff",
   72220 => x"ffffff",
   72221 => x"ffffff",
   72222 => x"ffffff",
   72223 => x"ffffff",
   72224 => x"ffffff",
   72225 => x"ffffff",
   72226 => x"ffffff",
   72227 => x"ffffff",
   72228 => x"ffffff",
   72229 => x"ffffff",
   72230 => x"ffffff",
   72231 => x"ffffff",
   72232 => x"ffffff",
   72233 => x"ffffff",
   72234 => x"ffffff",
   72235 => x"ffffff",
   72236 => x"ffffff",
   72237 => x"ffffff",
   72238 => x"ffffff",
   72239 => x"ffffff",
   72240 => x"ffffff",
   72241 => x"ffffff",
   72242 => x"ffffff",
   72243 => x"ffffff",
   72244 => x"ffffff",
   72245 => x"ffffff",
   72246 => x"ffffff",
   72247 => x"ffffff",
   72248 => x"ffffff",
   72249 => x"ffffff",
   72250 => x"ffffff",
   72251 => x"ffffff",
   72252 => x"ffffff",
   72253 => x"ffffff",
   72254 => x"ffffff",
   72255 => x"ffffff",
   72256 => x"ffffff",
   72257 => x"ffffff",
   72258 => x"ffffff",
   72259 => x"ffffff",
   72260 => x"ffffff",
   72261 => x"ffffff",
   72262 => x"ffffff",
   72263 => x"ffffff",
   72264 => x"ffffff",
   72265 => x"ffffff",
   72266 => x"ffffff",
   72267 => x"ffffff",
   72268 => x"ffffff",
   72269 => x"ffffff",
   72270 => x"ffffff",
   72271 => x"ffffff",
   72272 => x"ffffff",
   72273 => x"ffffff",
   72274 => x"ffffff",
   72275 => x"ffffff",
   72276 => x"ffffff",
   72277 => x"ffffff",
   72278 => x"ffffff",
   72279 => x"ffffff",
   72280 => x"ffffff",
   72281 => x"ffffff",
   72282 => x"ffffff",
   72283 => x"ffffff",
   72284 => x"ffffff",
   72285 => x"ffffff",
   72286 => x"ffffff",
   72287 => x"ffffff",
   72288 => x"ffffff",
   72289 => x"ffffff",
   72290 => x"ffffff",
   72291 => x"ffffff",
   72292 => x"ffffff",
   72293 => x"ffffff",
   72294 => x"ffffff",
   72295 => x"ffffff",
   72296 => x"ffffff",
   72297 => x"ffffff",
   72298 => x"ffffff",
   72299 => x"ffffff",
   72300 => x"ffffff",
   72301 => x"ffffff",
   72302 => x"ffffff",
   72303 => x"ffffff",
   72304 => x"ffffff",
   72305 => x"ffffff",
   72306 => x"ffffff",
   72307 => x"ffffff",
   72308 => x"ffffff",
   72309 => x"ffffff",
   72310 => x"ffffff",
   72311 => x"ffffff",
   72312 => x"ffffff",
   72313 => x"ffffff",
   72314 => x"ffffff",
   72315 => x"ffffff",
   72316 => x"ffffff",
   72317 => x"ffffff",
   72318 => x"ffffff",
   72319 => x"ffffff",
   72320 => x"ffffff",
   72321 => x"ffffff",
   72322 => x"ffffff",
   72323 => x"ffffff",
   72324 => x"ffffff",
   72325 => x"ffffff",
   72326 => x"ffffff",
   72327 => x"ffffff",
   72328 => x"ffffff",
   72329 => x"ffffff",
   72330 => x"ffffff",
   72331 => x"ffffff",
   72332 => x"ffffff",
   72333 => x"ffffff",
   72334 => x"ffffff",
   72335 => x"ffffff",
   72336 => x"ffffff",
   72337 => x"ffffff",
   72338 => x"ffffff",
   72339 => x"ffffff",
   72340 => x"ffffff",
   72341 => x"ffffff",
   72342 => x"ffffff",
   72343 => x"ffffff",
   72344 => x"ffffff",
   72345 => x"ffffff",
   72346 => x"ffffff",
   72347 => x"ffffff",
   72348 => x"ffffff",
   72349 => x"ffffff",
   72350 => x"ffffff",
   72351 => x"ffffff",
   72352 => x"ffffff",
   72353 => x"ffffff",
   72354 => x"ffffff",
   72355 => x"ffffff",
   72356 => x"ffffff",
   72357 => x"ffffff",
   72358 => x"ffffff",
   72359 => x"ffffff",
   72360 => x"ffffff",
   72361 => x"ffffff",
   72362 => x"ffffff",
   72363 => x"ffffff",
   72364 => x"ffffff",
   72365 => x"ffffff",
   72366 => x"ffffff",
   72367 => x"ffffff",
   72368 => x"ffffff",
   72369 => x"ffffff",
   72370 => x"ffffff",
   72371 => x"ffffff",
   72372 => x"ffffff",
   72373 => x"ffffff",
   72374 => x"ffffff",
   72375 => x"ffffff",
   72376 => x"ffffff",
   72377 => x"ffffff",
   72378 => x"ffffff",
   72379 => x"ffffff",
   72380 => x"ffffff",
   72381 => x"ffffff",
   72382 => x"ffffff",
   72383 => x"ffffff",
   72384 => x"ffffff",
   72385 => x"ffffff",
   72386 => x"ffffff",
   72387 => x"ffffff",
   72388 => x"ffffff",
   72389 => x"ffffff",
   72390 => x"ffffff",
   72391 => x"ffffff",
   72392 => x"ffffff",
   72393 => x"ffffff",
   72394 => x"ffffff",
   72395 => x"ffffff",
   72396 => x"ffffff",
   72397 => x"ffffff",
   72398 => x"ffffff",
   72399 => x"ffffff",
   72400 => x"ffffff",
   72401 => x"ffffff",
   72402 => x"ffffff",
   72403 => x"ffffff",
   72404 => x"ffffff",
   72405 => x"ffffff",
   72406 => x"ffffff",
   72407 => x"ffffff",
   72408 => x"ffffff",
   72409 => x"ffffff",
   72410 => x"ffffff",
   72411 => x"ffffff",
   72412 => x"ffffff",
   72413 => x"ffffff",
   72414 => x"ffffff",
   72415 => x"ffffff",
   72416 => x"ffffff",
   72417 => x"ffffff",
   72418 => x"ffffff",
   72419 => x"ffffff",
   72420 => x"ffffff",
   72421 => x"ffffff",
   72422 => x"ffffff",
   72423 => x"ffffff",
   72424 => x"ffffff",
   72425 => x"ffffff",
   72426 => x"ffffff",
   72427 => x"ffffff",
   72428 => x"ffffff",
   72429 => x"ffffff",
   72430 => x"ffffff",
   72431 => x"ffffff",
   72432 => x"ffffff",
   72433 => x"ffffff",
   72434 => x"ffffff",
   72435 => x"ffffff",
   72436 => x"ffffff",
   72437 => x"ffffff",
   72438 => x"ffffff",
   72439 => x"ffffff",
   72440 => x"ffffff",
   72441 => x"ffffff",
   72442 => x"ffffff",
   72443 => x"ffffff",
   72444 => x"ffffff",
   72445 => x"ffffff",
   72446 => x"ffffff",
   72447 => x"ffffff",
   72448 => x"ffffff",
   72449 => x"ffffff",
   72450 => x"ffffff",
   72451 => x"ffffff",
   72452 => x"ffffff",
   72453 => x"ffffff",
   72454 => x"ffffff",
   72455 => x"ffffff",
   72456 => x"ffffff",
   72457 => x"ffffff",
   72458 => x"ffffff",
   72459 => x"ffffff",
   72460 => x"ffffff",
   72461 => x"ffffff",
   72462 => x"ffffff",
   72463 => x"ffffff",
   72464 => x"ffffff",
   72465 => x"ffffff",
   72466 => x"ffffff",
   72467 => x"ffffff",
   72468 => x"ffffff",
   72469 => x"ffffff",
   72470 => x"ffffff",
   72471 => x"ffffff",
   72472 => x"ffffff",
   72473 => x"ffffff",
   72474 => x"ffffff",
   72475 => x"ffffff",
   72476 => x"ffffff",
   72477 => x"ffffff",
   72478 => x"ffffff",
   72479 => x"ffffff",
   72480 => x"ffffff",
   72481 => x"ffffff",
   72482 => x"ffffff",
   72483 => x"ffffff",
   72484 => x"ffffff",
   72485 => x"ffffff",
   72486 => x"ffffff",
   72487 => x"ffffff",
   72488 => x"ffffff",
   72489 => x"ffffff",
   72490 => x"ffffff",
   72491 => x"ffffff",
   72492 => x"ffffff",
   72493 => x"ffffff",
   72494 => x"ffffff",
   72495 => x"ffffff",
   72496 => x"ffffff",
   72497 => x"ffffff",
   72498 => x"ffffff",
   72499 => x"ffffff",
   72500 => x"ffffff",
   72501 => x"ffffff",
   72502 => x"ffffff",
   72503 => x"ffffff",
   72504 => x"ffffff",
   72505 => x"ffffff",
   72506 => x"ffffff",
   72507 => x"ffffff",
   72508 => x"ffffff",
   72509 => x"ffffff",
   72510 => x"ffffff",
   72511 => x"ffffff",
   72512 => x"ffffff",
   72513 => x"ffffff",
   72514 => x"ffffff",
   72515 => x"ffffff",
   72516 => x"ffffff",
   72517 => x"ffffff",
   72518 => x"ffffff",
   72519 => x"ffffff",
   72520 => x"ffffff",
   72521 => x"ffffff",
   72522 => x"ffffff",
   72523 => x"ffffff",
   72524 => x"ffffff",
   72525 => x"ffffff",
   72526 => x"ffffff",
   72527 => x"ffffff",
   72528 => x"ffffff",
   72529 => x"ffffff",
   72530 => x"ffffff",
   72531 => x"ffffff",
   72532 => x"ffffff",
   72533 => x"ffffff",
   72534 => x"ffffff",
   72535 => x"ffffff",
   72536 => x"ffffff",
   72537 => x"ffffff",
   72538 => x"ffffff",
   72539 => x"ffffff",
   72540 => x"ffffff",
   72541 => x"ffffff",
   72542 => x"ffffff",
   72543 => x"ffffff",
   72544 => x"ffffff",
   72545 => x"ffffff",
   72546 => x"ffffff",
   72547 => x"ffffff",
   72548 => x"ffffff",
   72549 => x"ffffff",
   72550 => x"ffffff",
   72551 => x"ffffff",
   72552 => x"ffffff",
   72553 => x"ffffff",
   72554 => x"ffffff",
   72555 => x"ffffff",
   72556 => x"ffffff",
   72557 => x"ffffff",
   72558 => x"ffffff",
   72559 => x"ffffff",
   72560 => x"ffffff",
   72561 => x"ffffff",
   72562 => x"ffffff",
   72563 => x"ffffff",
   72564 => x"ffffff",
   72565 => x"ffffff",
   72566 => x"ffffff",
   72567 => x"ffffff",
   72568 => x"ffffff",
   72569 => x"ffffff",
   72570 => x"ffffff",
   72571 => x"ffffff",
   72572 => x"ffffff",
   72573 => x"ffffff",
   72574 => x"ffffff",
   72575 => x"ffffff",
   72576 => x"ffffff",
   72577 => x"ffffff",
   72578 => x"ffffff",
   72579 => x"ffffff",
   72580 => x"ffffff",
   72581 => x"ffffff",
   72582 => x"ffffff",
   72583 => x"ffffff",
   72584 => x"ffffff",
   72585 => x"ffffff",
   72586 => x"ffffff",
   72587 => x"ffffff",
   72588 => x"ffffff",
   72589 => x"ffffff",
   72590 => x"ffffff",
   72591 => x"ffffff",
   72592 => x"ffffff",
   72593 => x"ffffff",
   72594 => x"ffffff",
   72595 => x"ffffff",
   72596 => x"ffffff",
   72597 => x"ffffff",
   72598 => x"ffffff",
   72599 => x"ffffff",
   72600 => x"ffffff",
   72601 => x"ffffff",
   72602 => x"ffffff",
   72603 => x"ffffff",
   72604 => x"ffffff",
   72605 => x"ffffff",
   72606 => x"ffffff",
   72607 => x"ffffff",
   72608 => x"ffffff",
   72609 => x"ffffff",
   72610 => x"ffffff",
   72611 => x"ffffff",
   72612 => x"ffffff",
   72613 => x"ffffff",
   72614 => x"ffffff",
   72615 => x"ffffff",
   72616 => x"ffffff",
   72617 => x"ffffff",
   72618 => x"ffffff",
   72619 => x"ffffff",
   72620 => x"ffffff",
   72621 => x"ffffff",
   72622 => x"ffffff",
   72623 => x"ffffff",
   72624 => x"ffffff",
   72625 => x"ffffff",
   72626 => x"ffffff",
   72627 => x"ffffff",
   72628 => x"ffffff",
   72629 => x"ffffff",
   72630 => x"ffffff",
   72631 => x"ffffff",
   72632 => x"ffffff",
   72633 => x"ffffff",
   72634 => x"ffffff",
   72635 => x"ffffff",
   72636 => x"ffffff",
   72637 => x"ffffff",
   72638 => x"ffffff",
   72639 => x"ffffff",
   72640 => x"ffffff",
   72641 => x"ffffff",
   72642 => x"ffffff",
   72643 => x"ffffff",
   72644 => x"ffffff",
   72645 => x"ffffff",
   72646 => x"ffffff",
   72647 => x"ffffff",
   72648 => x"ffffff",
   72649 => x"ffffff",
   72650 => x"ffffff",
   72651 => x"ffffff",
   72652 => x"ffffff",
   72653 => x"ffffff",
   72654 => x"ffffff",
   72655 => x"ffffff",
   72656 => x"ffffff",
   72657 => x"ffffff",
   72658 => x"ffffff",
   72659 => x"ffffff",
   72660 => x"ffffff",
   72661 => x"ffffff",
   72662 => x"ffffff",
   72663 => x"ffffff",
   72664 => x"ffffff",
   72665 => x"ffffff",
   72666 => x"ffffff",
   72667 => x"ffffff",
   72668 => x"ffffff",
   72669 => x"ffffff",
   72670 => x"ffffff",
   72671 => x"ffffff",
   72672 => x"ffffff",
   72673 => x"ffffff",
   72674 => x"ffffff",
   72675 => x"ffffff",
   72676 => x"ffffff",
   72677 => x"ffffff",
   72678 => x"ffffff",
   72679 => x"ffffff",
   72680 => x"ffffff",
   72681 => x"ffffff",
   72682 => x"ffffff",
   72683 => x"ffffff",
   72684 => x"ffffff",
   72685 => x"ffffff",
   72686 => x"ffffff",
   72687 => x"ffffff",
   72688 => x"ffffff",
   72689 => x"ffffff",
   72690 => x"ffffff",
   72691 => x"ffffff",
   72692 => x"ffffff",
   72693 => x"ffffff",
   72694 => x"ffffff",
   72695 => x"ffffff",
   72696 => x"ffffff",
   72697 => x"ffffff",
   72698 => x"ffffff",
   72699 => x"ffffff",
   72700 => x"ffffff",
   72701 => x"ffffff",
   72702 => x"ffffff",
   72703 => x"ffffff",
   72704 => x"ffffff",
   72705 => x"ffffff",
   72706 => x"ffffff",
   72707 => x"ffffff",
   72708 => x"ffffff",
   72709 => x"ffffff",
   72710 => x"ffffff",
   72711 => x"ffffff",
   72712 => x"ffffff",
   72713 => x"ffffff",
   72714 => x"ffffff",
   72715 => x"ffffff",
   72716 => x"ffffff",
   72717 => x"ffffff",
   72718 => x"ffffff",
   72719 => x"ffffff",
   72720 => x"ffffff",
   72721 => x"ffffff",
   72722 => x"ffffff",
   72723 => x"ffffff",
   72724 => x"ffffff",
   72725 => x"ffffff",
   72726 => x"ffffff",
   72727 => x"ffffff",
   72728 => x"ffffff",
   72729 => x"ffffff",
   72730 => x"ffffff",
   72731 => x"ffffff",
   72732 => x"ffffff",
   72733 => x"ffffff",
   72734 => x"ffffff",
   72735 => x"ffffff",
   72736 => x"ffffff",
   72737 => x"ffffff",
   72738 => x"ffffff",
   72739 => x"ffffff",
   72740 => x"ffffff",
   72741 => x"ffffff",
   72742 => x"ffffff",
   72743 => x"ffffff",
   72744 => x"ffffff",
   72745 => x"ffffff",
   72746 => x"ffffff",
   72747 => x"ffffff",
   72748 => x"ffffff",
   72749 => x"ffffff",
   72750 => x"ffffff",
   72751 => x"ffffff",
   72752 => x"ffffff",
   72753 => x"ffffff",
   72754 => x"ffffff",
   72755 => x"ffffff",
   72756 => x"ffffff",
   72757 => x"ffffff",
   72758 => x"ffffff",
   72759 => x"ffffff",
   72760 => x"ffffff",
   72761 => x"ffffff",
   72762 => x"ffffff",
   72763 => x"ffffff",
   72764 => x"ffffff",
   72765 => x"ffffff",
   72766 => x"ffffff",
   72767 => x"ffffff",
   72768 => x"ffffff",
   72769 => x"ffffff",
   72770 => x"ffffff",
   72771 => x"ffffff",
   72772 => x"ffffff",
   72773 => x"ffffff",
   72774 => x"ffffff",
   72775 => x"ffffff",
   72776 => x"ffffff",
   72777 => x"ffffff",
   72778 => x"ffffff",
   72779 => x"ffffff",
   72780 => x"ffffff",
   72781 => x"ffffff",
   72782 => x"ffffff",
   72783 => x"ffffff",
   72784 => x"ffffff",
   72785 => x"ffffff",
   72786 => x"ffffff",
   72787 => x"ffffff",
   72788 => x"ffffff",
   72789 => x"ffffff",
   72790 => x"ffffff",
   72791 => x"ffffff",
   72792 => x"ffffff",
   72793 => x"ffffff",
   72794 => x"ffffff",
   72795 => x"ffffff",
   72796 => x"ffffff",
   72797 => x"ffffff",
   72798 => x"ffffff",
   72799 => x"ffffff",
   72800 => x"ffffff",
   72801 => x"ffffff",
   72802 => x"ffffff",
   72803 => x"ffffff",
   72804 => x"ffffff",
   72805 => x"ffffff",
   72806 => x"ffffff",
   72807 => x"ffffff",
   72808 => x"ffffff",
   72809 => x"ffffff",
   72810 => x"ffffff",
   72811 => x"ffffff",
   72812 => x"ffffff",
   72813 => x"ffffff",
   72814 => x"ffffff",
   72815 => x"ffffff",
   72816 => x"ffffff",
   72817 => x"ffffff",
   72818 => x"ffffff",
   72819 => x"ffffff",
   72820 => x"ffffff",
   72821 => x"ffffff",
   72822 => x"ffffff",
   72823 => x"ffffff",
   72824 => x"ffffff",
   72825 => x"ffffff",
   72826 => x"ffffff",
   72827 => x"ffffff",
   72828 => x"ffffff",
   72829 => x"ffffff",
   72830 => x"ffffff",
   72831 => x"ffffff",
   72832 => x"ffffff",
   72833 => x"ffffff",
   72834 => x"ffffff",
   72835 => x"ffffff",
   72836 => x"ffffff",
   72837 => x"ffffff",
   72838 => x"ffffff",
   72839 => x"ffffff",
   72840 => x"ffffff",
   72841 => x"ffffff",
   72842 => x"ffffff",
   72843 => x"ffffff",
   72844 => x"ffffff",
   72845 => x"ffffff",
   72846 => x"ffffff",
   72847 => x"ffffff",
   72848 => x"ffffff",
   72849 => x"ffffff",
   72850 => x"ffffff",
   72851 => x"ffffff",
   72852 => x"ffffff",
   72853 => x"ffffff",
   72854 => x"ffffff",
   72855 => x"ffffff",
   72856 => x"ffffff",
   72857 => x"ffffff",
   72858 => x"ffffff",
   72859 => x"ffffff",
   72860 => x"ffffff",
   72861 => x"ffffff",
   72862 => x"ffffff",
   72863 => x"ffffff",
   72864 => x"ffffff",
   72865 => x"ffffff",
   72866 => x"ffffff",
   72867 => x"ffffff",
   72868 => x"ffffff",
   72869 => x"ffffff",
   72870 => x"ffffff",
   72871 => x"ffffff",
   72872 => x"ffffff",
   72873 => x"ffffff",
   72874 => x"ffffff",
   72875 => x"ffffff",
   72876 => x"ffffff",
   72877 => x"ffffff",
   72878 => x"ffffff",
   72879 => x"ffffff",
   72880 => x"ffffff",
   72881 => x"ffffff",
   72882 => x"ffffff",
   72883 => x"ffffff",
   72884 => x"ffffff",
   72885 => x"ffffff",
   72886 => x"ffffff",
   72887 => x"ffffff",
   72888 => x"ffffff",
   72889 => x"ffffff",
   72890 => x"ffffff",
   72891 => x"ffffff",
   72892 => x"ffffff",
   72893 => x"ffffff",
   72894 => x"ffffff",
   72895 => x"ffffff",
   72896 => x"ffffff",
   72897 => x"ffffff",
   72898 => x"ffffff",
   72899 => x"ffffff",
   72900 => x"ffffff",
   72901 => x"ffffff",
   72902 => x"ffffff",
   72903 => x"ffffff",
   72904 => x"ffffff",
   72905 => x"ffffff",
   72906 => x"ffffff",
   72907 => x"ffffff",
   72908 => x"ffffff",
   72909 => x"ffffff",
   72910 => x"ffffff",
   72911 => x"ffffff",
   72912 => x"ffffff",
   72913 => x"ffffff",
   72914 => x"ffffff",
   72915 => x"ffffff",
   72916 => x"ffffff",
   72917 => x"ffffff",
   72918 => x"ffffff",
   72919 => x"ffffff",
   72920 => x"ffffff",
   72921 => x"ffffff",
   72922 => x"ffffff",
   72923 => x"ffffff",
   72924 => x"ffffff",
   72925 => x"ffffff",
   72926 => x"ffffff",
   72927 => x"ffffff",
   72928 => x"ffffff",
   72929 => x"ffffff",
   72930 => x"ffffff",
   72931 => x"ffffff",
   72932 => x"ffffff",
   72933 => x"ffffff",
   72934 => x"ffffff",
   72935 => x"ffffff",
   72936 => x"ffffff",
   72937 => x"ffffff",
   72938 => x"ffffff",
   72939 => x"ffffff",
   72940 => x"ffffff",
   72941 => x"ffffff",
   72942 => x"ffffff",
   72943 => x"ffffff",
   72944 => x"ffffff",
   72945 => x"ffffff",
   72946 => x"ffffff",
   72947 => x"ffffff",
   72948 => x"ffffff",
   72949 => x"ffffff",
   72950 => x"ffffff",
   72951 => x"ffffff",
   72952 => x"ffffff",
   72953 => x"ffffff",
   72954 => x"ffffff",
   72955 => x"ffffff",
   72956 => x"ffffff",
   72957 => x"ffffff",
   72958 => x"ffffff",
   72959 => x"ffffff",
   72960 => x"ffffff",
   72961 => x"ffffff",
   72962 => x"ffffff",
   72963 => x"ffffff",
   72964 => x"ffffff",
   72965 => x"ffffff",
   72966 => x"ffffff",
   72967 => x"ffffff",
   72968 => x"ffffff",
   72969 => x"ffffff",
   72970 => x"ffffff",
   72971 => x"ffffff",
   72972 => x"ffffff",
   72973 => x"ffffff",
   72974 => x"ffffff",
   72975 => x"ffffff",
   72976 => x"ffffff",
   72977 => x"ffffff",
   72978 => x"ffffff",
   72979 => x"ffffff",
   72980 => x"ffffff",
   72981 => x"ffffff",
   72982 => x"ffffff",
   72983 => x"ffffff",
   72984 => x"ffffff",
   72985 => x"ffffff",
   72986 => x"ffffff",
   72987 => x"ffffff",
   72988 => x"ffffff",
   72989 => x"ffffff",
   72990 => x"ffffff",
   72991 => x"ffffff",
   72992 => x"ffffff",
   72993 => x"ffffff",
   72994 => x"ffffff",
   72995 => x"ffffff",
   72996 => x"ffffff",
   72997 => x"ffffff",
   72998 => x"ffffff",
   72999 => x"ffffff",
   73000 => x"ffffff",
   73001 => x"ffffff",
   73002 => x"ffffff",
   73003 => x"ffffff",
   73004 => x"ffffff",
   73005 => x"ffffff",
   73006 => x"ffffff",
   73007 => x"ffffff",
   73008 => x"ffffff",
   73009 => x"ffffff",
   73010 => x"ffffff",
   73011 => x"ffffff",
   73012 => x"ffffff",
   73013 => x"ffffff",
   73014 => x"ffffff",
   73015 => x"ffffff",
   73016 => x"ffffff",
   73017 => x"ffffff",
   73018 => x"ffffff",
   73019 => x"ffffff",
   73020 => x"ffffff",
   73021 => x"ffffff",
   73022 => x"ffffff",
   73023 => x"ffffff",
   73024 => x"ffffff",
   73025 => x"ffffff",
   73026 => x"ffffff",
   73027 => x"ffffff",
   73028 => x"ffffff",
   73029 => x"ffffff",
   73030 => x"ffffff",
   73031 => x"ffffff",
   73032 => x"ffffff",
   73033 => x"ffffff",
   73034 => x"ffffff",
   73035 => x"ffffff",
   73036 => x"ffffff",
   73037 => x"ffffff",
   73038 => x"ffffff",
   73039 => x"ffffff",
   73040 => x"ffffff",
   73041 => x"ffffff",
   73042 => x"ffffff",
   73043 => x"ffffff",
   73044 => x"ffffff",
   73045 => x"ffffff",
   73046 => x"ffffff",
   73047 => x"ffffff",
   73048 => x"ffffff",
   73049 => x"ffffff",
   73050 => x"ffffff",
   73051 => x"ffffff",
   73052 => x"ffffff",
   73053 => x"ffffff",
   73054 => x"ffffff",
   73055 => x"ffffff",
   73056 => x"ffffff",
   73057 => x"ffffff",
   73058 => x"ffffff",
   73059 => x"ffffff",
   73060 => x"ffffff",
   73061 => x"ffffff",
   73062 => x"ffffff",
   73063 => x"ffffff",
   73064 => x"ffffff",
   73065 => x"ffffff",
   73066 => x"ffffff",
   73067 => x"ffffff",
   73068 => x"ffffff",
   73069 => x"ffffff",
   73070 => x"ffffff",
   73071 => x"ffffff",
   73072 => x"ffffff",
   73073 => x"ffffff",
   73074 => x"ffffff",
   73075 => x"ffffff",
   73076 => x"ffffff",
   73077 => x"ffffff",
   73078 => x"ffffff",
   73079 => x"ffffff",
   73080 => x"ffffff",
   73081 => x"ffffff",
   73082 => x"ffffff",
   73083 => x"ffffff",
   73084 => x"ffffff",
   73085 => x"ffffff",
   73086 => x"ffffff",
   73087 => x"ffffff",
   73088 => x"ffffff",
   73089 => x"ffffff",
   73090 => x"ffffff",
   73091 => x"ffffff",
   73092 => x"ffffff",
   73093 => x"ffffff",
   73094 => x"ffffff",
   73095 => x"ffffff",
   73096 => x"ffffff",
   73097 => x"ffffff",
   73098 => x"ffffff",
   73099 => x"ffffff",
   73100 => x"ffffff",
   73101 => x"ffffff",
   73102 => x"ffffff",
   73103 => x"ffffff",
   73104 => x"ffffff",
   73105 => x"ffffff",
   73106 => x"ffffff",
   73107 => x"ffffff",
   73108 => x"ffffff",
   73109 => x"ffffff",
   73110 => x"ffffff",
   73111 => x"ffffff",
   73112 => x"ffffff",
   73113 => x"ffffff",
   73114 => x"ffffff",
   73115 => x"ffffff",
   73116 => x"ffffff",
   73117 => x"ffffff",
   73118 => x"ffffff",
   73119 => x"ffffff",
   73120 => x"ffffff",
   73121 => x"ffffff",
   73122 => x"ffffff",
   73123 => x"ffffff",
   73124 => x"ffffff",
   73125 => x"ffffff",
   73126 => x"ffffff",
   73127 => x"ffffff",
   73128 => x"ffffff",
   73129 => x"ffffff",
   73130 => x"ffffff",
   73131 => x"ffffff",
   73132 => x"ffffff",
   73133 => x"ffffff",
   73134 => x"ffffff",
   73135 => x"ffffff",
   73136 => x"ffffff",
   73137 => x"ffffff",
   73138 => x"ffffff",
   73139 => x"ffffff",
   73140 => x"ffffff",
   73141 => x"ffffff",
   73142 => x"ffffff",
   73143 => x"ffffff",
   73144 => x"ffffff",
   73145 => x"ffffff",
   73146 => x"ffffff",
   73147 => x"ffffff",
   73148 => x"ffffff",
   73149 => x"ffffff",
   73150 => x"ffffff",
   73151 => x"ffffff",
   73152 => x"ffffff",
   73153 => x"ffffff",
   73154 => x"ffffff",
   73155 => x"ffffff",
   73156 => x"ffffff",
   73157 => x"ffffff",
   73158 => x"ffffff",
   73159 => x"ffffff",
   73160 => x"ffffff",
   73161 => x"ffffff",
   73162 => x"ffffff",
   73163 => x"ffffff",
   73164 => x"ffffff",
   73165 => x"ffffff",
   73166 => x"ffffff",
   73167 => x"ffffff",
   73168 => x"ffffff",
   73169 => x"ffffff",
   73170 => x"ffffff",
   73171 => x"ffffff",
   73172 => x"ffffff",
   73173 => x"ffffff",
   73174 => x"ffffff",
   73175 => x"ffffff",
   73176 => x"ffffff",
   73177 => x"ffffff",
   73178 => x"ffffff",
   73179 => x"ffffff",
   73180 => x"ffffff",
   73181 => x"ffffff",
   73182 => x"ffffff",
   73183 => x"ffffff",
   73184 => x"ffffff",
   73185 => x"ffffff",
   73186 => x"ffffff",
   73187 => x"ffffff",
   73188 => x"ffffff",
   73189 => x"ffffff",
   73190 => x"ffffff",
   73191 => x"ffffff",
   73192 => x"ffffff",
   73193 => x"ffffff",
   73194 => x"ffffff",
   73195 => x"ffffff",
   73196 => x"ffffff",
   73197 => x"ffffff",
   73198 => x"ffffff",
   73199 => x"ffffff",
   73200 => x"ffffff",
   73201 => x"ffffff",
   73202 => x"ffffff",
   73203 => x"ffffff",
   73204 => x"ffffff",
   73205 => x"ffffff",
   73206 => x"ffffff",
   73207 => x"ffffff",
   73208 => x"ffffff",
   73209 => x"ffffff",
   73210 => x"ffffff",
   73211 => x"ffffff",
   73212 => x"ffffff",
   73213 => x"ffffff",
   73214 => x"ffffff",
   73215 => x"ffffff",
   73216 => x"ffffff",
   73217 => x"ffffff",
   73218 => x"ffffff",
   73219 => x"ffffff",
   73220 => x"ffffff",
   73221 => x"ffffff",
   73222 => x"ffffff",
   73223 => x"ffffff",
   73224 => x"ffffff",
   73225 => x"ffffff",
   73226 => x"ffffff",
   73227 => x"ffffff",
   73228 => x"ffffff",
   73229 => x"ffffff",
   73230 => x"ffffff",
   73231 => x"ffffff",
   73232 => x"ffffff",
   73233 => x"ffffff",
   73234 => x"ffffff",
   73235 => x"ffffff",
   73236 => x"ffffff",
   73237 => x"ffffff",
   73238 => x"ffffff",
   73239 => x"ffffff",
   73240 => x"ffffff",
   73241 => x"ffffff",
   73242 => x"ffffff",
   73243 => x"ffffff",
   73244 => x"ffffff",
   73245 => x"ffffff",
   73246 => x"ffffff",
   73247 => x"ffffff",
   73248 => x"ffffff",
   73249 => x"ffffff",
   73250 => x"ffffff",
   73251 => x"ffffff",
   73252 => x"ffffff",
   73253 => x"ffffff",
   73254 => x"ffffff",
   73255 => x"ffffff",
   73256 => x"ffffff",
   73257 => x"ffffff",
   73258 => x"ffffff",
   73259 => x"ffffff",
   73260 => x"ffffff",
   73261 => x"ffffff",
   73262 => x"ffffff",
   73263 => x"ffffff",
   73264 => x"ffffff",
   73265 => x"ffffff",
   73266 => x"ffffff",
   73267 => x"ffffff",
   73268 => x"ffffff",
   73269 => x"ffffff",
   73270 => x"ffffff",
   73271 => x"ffffff",
   73272 => x"ffffff",
   73273 => x"ffffff",
   73274 => x"ffffff",
   73275 => x"ffffff",
   73276 => x"ffffff",
   73277 => x"ffffff",
   73278 => x"ffffff",
   73279 => x"ffffff",
   73280 => x"ffffff",
   73281 => x"ffffff",
   73282 => x"ffffff",
   73283 => x"ffffff",
   73284 => x"ffffff",
   73285 => x"ffffff",
   73286 => x"ffffff",
   73287 => x"ffffff",
   73288 => x"ffffff",
   73289 => x"ffffff",
   73290 => x"ffffff",
   73291 => x"ffffff",
   73292 => x"ffffff",
   73293 => x"ffffff",
   73294 => x"ffffff",
   73295 => x"ffffff",
   73296 => x"ffffff",
   73297 => x"ffffff",
   73298 => x"ffffff",
   73299 => x"ffffff",
   73300 => x"ffffff",
   73301 => x"ffffff",
   73302 => x"ffffff",
   73303 => x"ffffff",
   73304 => x"ffffff",
   73305 => x"ffffff",
   73306 => x"ffffff",
   73307 => x"ffffff",
   73308 => x"ffffff",
   73309 => x"ffffff",
   73310 => x"ffffff",
   73311 => x"ffffff",
   73312 => x"ffffff",
   73313 => x"ffffff",
   73314 => x"ffffff",
   73315 => x"ffffff",
   73316 => x"ffffff",
   73317 => x"ffffff",
   73318 => x"ffffff",
   73319 => x"ffffff",
   73320 => x"ffffff",
   73321 => x"ffffff",
   73322 => x"ffffff",
   73323 => x"ffffff",
   73324 => x"ffffff",
   73325 => x"ffffff",
   73326 => x"ffffff",
   73327 => x"ffffff",
   73328 => x"ffffff",
   73329 => x"ffffff",
   73330 => x"ffffff",
   73331 => x"ffffff",
   73332 => x"ffffff",
   73333 => x"ffffff",
   73334 => x"ffffff",
   73335 => x"ffffff",
   73336 => x"ffffff",
   73337 => x"ffffff",
   73338 => x"ffffff",
   73339 => x"ffffff",
   73340 => x"ffffff",
   73341 => x"ffffff",
   73342 => x"ffffff",
   73343 => x"ffffff",
   73344 => x"ffffff",
   73345 => x"ffffff",
   73346 => x"ffffff",
   73347 => x"ffffff",
   73348 => x"ffffff",
   73349 => x"ffffff",
   73350 => x"ffffff",
   73351 => x"ffffff",
   73352 => x"ffffff",
   73353 => x"ffffff",
   73354 => x"ffffff",
   73355 => x"ffffff",
   73356 => x"ffffff",
   73357 => x"ffffff",
   73358 => x"ffffff",
   73359 => x"ffffff",
   73360 => x"ffffff",
   73361 => x"ffffff",
   73362 => x"ffffff",
   73363 => x"ffffff",
   73364 => x"ffffff",
   73365 => x"ffffff",
   73366 => x"ffffff",
   73367 => x"ffffff",
   73368 => x"ffffff",
   73369 => x"ffffff",
   73370 => x"ffffff",
   73371 => x"ffffff",
   73372 => x"ffffff",
   73373 => x"ffffff",
   73374 => x"ffffff",
   73375 => x"ffffff",
   73376 => x"ffffff",
   73377 => x"ffffff",
   73378 => x"ffffff",
   73379 => x"ffffff",
   73380 => x"ffffff",
   73381 => x"ffffff",
   73382 => x"ffffff",
   73383 => x"ffffff",
   73384 => x"ffffff",
   73385 => x"ffffff",
   73386 => x"ffffff",
   73387 => x"ffffff",
   73388 => x"ffffff",
   73389 => x"ffffff",
   73390 => x"ffffff",
   73391 => x"ffffff",
   73392 => x"ffffff",
   73393 => x"ffffff",
   73394 => x"ffffff",
   73395 => x"ffffff",
   73396 => x"ffffff",
   73397 => x"ffffff",
   73398 => x"ffffff",
   73399 => x"ffffff",
   73400 => x"ffffff",
   73401 => x"ffffff",
   73402 => x"ffffff",
   73403 => x"ffffff",
   73404 => x"ffffff",
   73405 => x"ffffff",
   73406 => x"ffffff",
   73407 => x"ffffff",
   73408 => x"ffffff",
   73409 => x"ffffff",
   73410 => x"ffffff",
   73411 => x"ffffff",
   73412 => x"ffffff",
   73413 => x"ffffff",
   73414 => x"ffffff",
   73415 => x"ffffff",
   73416 => x"ffffff",
   73417 => x"ffffff",
   73418 => x"ffffff",
   73419 => x"ffffff",
   73420 => x"ffffff",
   73421 => x"ffffff",
   73422 => x"ffffff",
   73423 => x"ffffff",
   73424 => x"ffffff",
   73425 => x"ffffff",
   73426 => x"ffffff",
   73427 => x"ffffff",
   73428 => x"ffffff",
   73429 => x"ffffff",
   73430 => x"ffffff",
   73431 => x"ffffff",
   73432 => x"ffffff",
   73433 => x"ffffff",
   73434 => x"ffffff",
   73435 => x"ffffff",
   73436 => x"ffffff",
   73437 => x"ffffff",
   73438 => x"ffffff",
   73439 => x"ffffff",
   73440 => x"ffffff",
   73441 => x"ffffff",
   73442 => x"ffffff",
   73443 => x"ffffff",
   73444 => x"ffffff",
   73445 => x"ffffff",
   73446 => x"ffffff",
   73447 => x"ffffff",
   73448 => x"ffffff",
   73449 => x"ffffff",
   73450 => x"ffffff",
   73451 => x"ffffff",
   73452 => x"ffffff",
   73453 => x"ffffff",
   73454 => x"ffffff",
   73455 => x"ffffff",
   73456 => x"ffffff",
   73457 => x"ffffff",
   73458 => x"ffffff",
   73459 => x"ffffff",
   73460 => x"ffffff",
   73461 => x"ffffff",
   73462 => x"ffffff",
   73463 => x"ffffff",
   73464 => x"ffffff",
   73465 => x"ffffff",
   73466 => x"ffffff",
   73467 => x"ffffff",
   73468 => x"ffffff",
   73469 => x"ffffff",
   73470 => x"ffffff",
   73471 => x"ffffff",
   73472 => x"ffffff",
   73473 => x"ffffff",
   73474 => x"ffffff",
   73475 => x"ffffff",
   73476 => x"ffffff",
   73477 => x"ffffff",
   73478 => x"ffffff",
   73479 => x"ffffff",
   73480 => x"ffffff",
   73481 => x"ffffff",
   73482 => x"ffffff",
   73483 => x"ffffff",
   73484 => x"ffffff",
   73485 => x"ffffff",
   73486 => x"ffffff",
   73487 => x"ffffff",
   73488 => x"ffffff",
   73489 => x"ffffff",
   73490 => x"ffffff",
   73491 => x"ffffff",
   73492 => x"ffffff",
   73493 => x"ffffff",
   73494 => x"ffffff",
   73495 => x"ffffff",
   73496 => x"ffffff",
   73497 => x"ffffff",
   73498 => x"ffffff",
   73499 => x"ffffff",
   73500 => x"ffffff",
   73501 => x"ffffff",
   73502 => x"ffffff",
   73503 => x"ffffff",
   73504 => x"ffffff",
   73505 => x"ffffff",
   73506 => x"ffffff",
   73507 => x"ffffff",
   73508 => x"ffffff",
   73509 => x"ffffff",
   73510 => x"ffffff",
   73511 => x"ffffff",
   73512 => x"ffffff",
   73513 => x"ffffff",
   73514 => x"ffffff",
   73515 => x"ffffff",
   73516 => x"ffffff",
   73517 => x"ffffff",
   73518 => x"ffffff",
   73519 => x"ffffff",
   73520 => x"ffffff",
   73521 => x"ffffff",
   73522 => x"ffffff",
   73523 => x"ffffff",
   73524 => x"ffffff",
   73525 => x"ffffff",
   73526 => x"ffffff",
   73527 => x"ffffff",
   73528 => x"ffffff",
   73529 => x"ffffff",
   73530 => x"ffffff",
   73531 => x"ffffff",
   73532 => x"ffffff",
   73533 => x"ffffff",
   73534 => x"ffffff",
   73535 => x"ffffff",
   73536 => x"ffffff",
   73537 => x"ffffff",
   73538 => x"ffffff",
   73539 => x"ffffff",
   73540 => x"ffffff",
   73541 => x"ffffff",
   73542 => x"ffffff",
   73543 => x"ffffff",
   73544 => x"ffffff",
   73545 => x"ffffff",
   73546 => x"ffffff",
   73547 => x"ffffff",
   73548 => x"ffffff",
   73549 => x"ffffff",
   73550 => x"ffffff",
   73551 => x"ffffff",
   73552 => x"ffffff",
   73553 => x"ffffff",
   73554 => x"ffffff",
   73555 => x"ffffff",
   73556 => x"ffffff",
   73557 => x"ffffff",
   73558 => x"ffffff",
   73559 => x"ffffff",
   73560 => x"ffffff",
   73561 => x"ffffff",
   73562 => x"ffffff",
   73563 => x"ffffff",
   73564 => x"ffffff",
   73565 => x"ffffff",
   73566 => x"ffffff",
   73567 => x"ffffff",
   73568 => x"ffffff",
   73569 => x"ffffff",
   73570 => x"ffffff",
   73571 => x"ffffff",
   73572 => x"ffffff",
   73573 => x"ffffff",
   73574 => x"ffffff",
   73575 => x"ffffff",
   73576 => x"ffffff",
   73577 => x"ffffff",
   73578 => x"ffffff",
   73579 => x"ffffff",
   73580 => x"ffffff",
   73581 => x"ffffff",
   73582 => x"ffffff",
   73583 => x"ffffff",
   73584 => x"ffffff",
   73585 => x"ffffff",
   73586 => x"ffffff",
   73587 => x"ffffff",
   73588 => x"ffffff",
   73589 => x"ffffff",
   73590 => x"ffffff",
   73591 => x"ffffff",
   73592 => x"ffffff",
   73593 => x"ffffff",
   73594 => x"ffffff",
   73595 => x"ffffff",
   73596 => x"ffffff",
   73597 => x"ffffff",
   73598 => x"ffffff",
   73599 => x"ffffff",
   73600 => x"ffffff",
   73601 => x"ffffff",
   73602 => x"ffffff",
   73603 => x"ffffff",
   73604 => x"ffffff",
   73605 => x"ffffff",
   73606 => x"ffffff",
   73607 => x"ffffff",
   73608 => x"ffffff",
   73609 => x"ffffff",
   73610 => x"ffffff",
   73611 => x"ffffff",
   73612 => x"ffffff",
   73613 => x"ffffff",
   73614 => x"ffffff",
   73615 => x"ffffff",
   73616 => x"ffffff",
   73617 => x"ffffff",
   73618 => x"ffffff",
   73619 => x"ffffff",
   73620 => x"ffffff",
   73621 => x"ffffff",
   73622 => x"ffffff",
   73623 => x"ffffff",
   73624 => x"ffffff",
   73625 => x"ffffff",
   73626 => x"ffffff",
   73627 => x"ffffff",
   73628 => x"ffffff",
   73629 => x"ffffff",
   73630 => x"ffffff",
   73631 => x"ffffff",
   73632 => x"ffffff",
   73633 => x"ffffff",
   73634 => x"ffffff",
   73635 => x"ffffff",
   73636 => x"ffffff",
   73637 => x"ffffff",
   73638 => x"ffffff",
   73639 => x"ffffff",
   73640 => x"ffffff",
   73641 => x"ffffff",
   73642 => x"ffffff",
   73643 => x"ffffff",
   73644 => x"ffffff",
   73645 => x"ffffff",
   73646 => x"ffffff",
   73647 => x"ffffff",
   73648 => x"ffffff",
   73649 => x"ffffff",
   73650 => x"ffffff",
   73651 => x"ffffff",
   73652 => x"ffffff",
   73653 => x"ffffff",
   73654 => x"ffffff",
   73655 => x"ffffff",
   73656 => x"ffffff",
   73657 => x"ffffff",
   73658 => x"ffffff",
   73659 => x"ffffff",
   73660 => x"ffffff",
   73661 => x"ffffff",
   73662 => x"ffffff",
   73663 => x"ffffff",
   73664 => x"ffffff",
   73665 => x"ffffff",
   73666 => x"ffffff",
   73667 => x"ffffff",
   73668 => x"ffffff",
   73669 => x"ffffff",
   73670 => x"ffffff",
   73671 => x"ffffff",
   73672 => x"ffffff",
   73673 => x"ffffff",
   73674 => x"ffffff",
   73675 => x"ffffff",
   73676 => x"ffffff",
   73677 => x"ffffff",
   73678 => x"ffffff",
   73679 => x"ffffff",
   73680 => x"ffffff",
   73681 => x"ffffff",
   73682 => x"ffffff",
   73683 => x"ffffff",
   73684 => x"ffffff",
   73685 => x"ffffff",
   73686 => x"ffffff",
   73687 => x"ffffff",
   73688 => x"ffffff",
   73689 => x"ffffff",
   73690 => x"ffffff",
   73691 => x"ffffff",
   73692 => x"ffffff",
   73693 => x"ffffff",
   73694 => x"ffffff",
   73695 => x"ffffff",
   73696 => x"ffffff",
   73697 => x"ffffff",
   73698 => x"ffffff",
   73699 => x"ffffff",
   73700 => x"ffffff",
   73701 => x"ffffff",
   73702 => x"ffffff",
   73703 => x"ffffff",
   73704 => x"ffffff",
   73705 => x"ffffff",
   73706 => x"ffffff",
   73707 => x"ffffff",
   73708 => x"ffffff",
   73709 => x"ffffff",
   73710 => x"ffffff",
   73711 => x"ffffff",
   73712 => x"ffffff",
   73713 => x"ffffff",
   73714 => x"ffffff",
   73715 => x"ffffff",
   73716 => x"ffffff",
   73717 => x"ffffff",
   73718 => x"ffffff",
   73719 => x"ffffff",
   73720 => x"ffffff",
   73721 => x"ffffff",
   73722 => x"ffffff",
   73723 => x"ffffff",
   73724 => x"ffffff",
   73725 => x"ffffff",
   73726 => x"ffffff",
   73727 => x"ffffff",
   73728 => x"ffffff",
   73729 => x"ffffff",
   73730 => x"ffffff",
   73731 => x"ffffff",
   73732 => x"ffffff",
   73733 => x"ffffff",
   73734 => x"ffffff",
   73735 => x"ffffff",
   73736 => x"ffffff",
   73737 => x"ffffff",
   73738 => x"ffffff",
   73739 => x"ffffff",
   73740 => x"ffffff",
   73741 => x"ffffff",
   73742 => x"ffffff",
   73743 => x"ffffff",
   73744 => x"ffffff",
   73745 => x"ffffff",
   73746 => x"ffffff",
   73747 => x"ffffff",
   73748 => x"ffffff",
   73749 => x"ffffff",
   73750 => x"ffffff",
   73751 => x"ffffff",
   73752 => x"ffffff",
   73753 => x"ffffff",
   73754 => x"ffffff",
   73755 => x"ffffff",
   73756 => x"ffffff",
   73757 => x"ffffff",
   73758 => x"ffffff",
   73759 => x"ffffff",
   73760 => x"ffffff",
   73761 => x"ffffff",
   73762 => x"ffffff",
   73763 => x"ffffff",
   73764 => x"ffffff",
   73765 => x"ffffff",
   73766 => x"ffffff",
   73767 => x"ffffff",
   73768 => x"ffffff",
   73769 => x"ffffff",
   73770 => x"ffffff",
   73771 => x"ffffff",
   73772 => x"ffffff",
   73773 => x"ffffff",
   73774 => x"ffffff",
   73775 => x"ffffff",
   73776 => x"ffffff",
   73777 => x"ffffff",
   73778 => x"ffffff",
   73779 => x"ffffff",
   73780 => x"ffffff",
   73781 => x"ffffff",
   73782 => x"ffffff",
   73783 => x"ffffff",
   73784 => x"ffffff",
   73785 => x"ffffff",
   73786 => x"ffffff",
   73787 => x"ffffff",
   73788 => x"ffffff",
   73789 => x"ffffff",
   73790 => x"ffffff",
   73791 => x"ffffff",
   73792 => x"ffffff",
   73793 => x"ffffff",
   73794 => x"ffffff",
   73795 => x"ffffff",
   73796 => x"ffffff",
   73797 => x"ffffff",
   73798 => x"ffffff",
   73799 => x"ffffff",
   73800 => x"ffffff",
   73801 => x"ffffff",
   73802 => x"ffffff",
   73803 => x"ffffff",
   73804 => x"ffffff",
   73805 => x"ffffff",
   73806 => x"ffffff",
   73807 => x"ffffff",
   73808 => x"ffffff",
   73809 => x"ffffff",
   73810 => x"ffffff",
   73811 => x"ffffff",
   73812 => x"ffffff",
   73813 => x"ffffff",
   73814 => x"ffffff",
   73815 => x"ffffff",
   73816 => x"ffffff",
   73817 => x"ffffff",
   73818 => x"ffffff",
   73819 => x"ffffff",
   73820 => x"ffffff",
   73821 => x"ffffff",
   73822 => x"ffffff",
   73823 => x"ffffff",
   73824 => x"ffffff",
   73825 => x"ffffff",
   73826 => x"ffffff",
   73827 => x"ffffff",
   73828 => x"ffffff",
   73829 => x"ffffff",
   73830 => x"ffffff",
   73831 => x"ffffff",
   73832 => x"ffffff",
   73833 => x"ffffff",
   73834 => x"ffffff",
   73835 => x"ffffff",
   73836 => x"ffffff",
   73837 => x"ffffff",
   73838 => x"ffffff",
   73839 => x"ffffff",
   73840 => x"ffffff",
   73841 => x"ffffff",
   73842 => x"ffffff",
   73843 => x"ffffff",
   73844 => x"ffffff",
   73845 => x"ffffff",
   73846 => x"ffffff",
   73847 => x"ffffff",
   73848 => x"ffffff",
   73849 => x"ffffff",
   73850 => x"ffffff",
   73851 => x"ffffff",
   73852 => x"ffffff",
   73853 => x"ffffff",
   73854 => x"ffffff",
   73855 => x"ffffff",
   73856 => x"ffffff",
   73857 => x"ffffff",
   73858 => x"ffffff",
   73859 => x"ffffff",
   73860 => x"ffffff",
   73861 => x"ffffff",
   73862 => x"ffffff",
   73863 => x"ffffff",
   73864 => x"ffffff",
   73865 => x"ffffff",
   73866 => x"ffffff",
   73867 => x"ffffff",
   73868 => x"ffffff",
   73869 => x"ffffff",
   73870 => x"ffffff",
   73871 => x"ffffff",
   73872 => x"ffffff",
   73873 => x"ffffff",
   73874 => x"ffffff",
   73875 => x"ffffff",
   73876 => x"ffffff",
   73877 => x"ffffff",
   73878 => x"ffffff",
   73879 => x"ffffff",
   73880 => x"ffffff",
   73881 => x"ffffff",
   73882 => x"ffffff",
   73883 => x"ffffff",
   73884 => x"ffffff",
   73885 => x"ffffff",
   73886 => x"ffffff",
   73887 => x"ffffff",
   73888 => x"ffffff",
   73889 => x"ffffff",
   73890 => x"ffffff",
   73891 => x"ffffff",
   73892 => x"ffffff",
   73893 => x"ffffff",
   73894 => x"ffffff",
   73895 => x"ffffff",
   73896 => x"ffffff",
   73897 => x"ffffff",
   73898 => x"ffffff",
   73899 => x"ffffff",
   73900 => x"ffffff",
   73901 => x"ffffff",
   73902 => x"ffffff",
   73903 => x"ffffff",
   73904 => x"ffffff",
   73905 => x"ffffff",
   73906 => x"ffffff",
   73907 => x"ffffff",
   73908 => x"ffffff",
   73909 => x"ffffff",
   73910 => x"ffffff",
   73911 => x"ffffff",
   73912 => x"ffffff",
   73913 => x"ffffff",
   73914 => x"ffffff",
   73915 => x"ffffff",
   73916 => x"ffffff",
   73917 => x"ffffff",
   73918 => x"ffffff",
   73919 => x"ffffff",
   73920 => x"ffffff",
   73921 => x"ffffff",
   73922 => x"ffffff",
   73923 => x"ffffff",
   73924 => x"ffffff",
   73925 => x"ffffff",
   73926 => x"ffffff",
   73927 => x"ffffff",
   73928 => x"ffffff",
   73929 => x"ffffff",
   73930 => x"ffffff",
   73931 => x"ffffff",
   73932 => x"ffffff",
   73933 => x"ffffff",
   73934 => x"ffffff",
   73935 => x"ffffff",
   73936 => x"ffffff",
   73937 => x"ffffff",
   73938 => x"ffffff",
   73939 => x"ffffff",
   73940 => x"ffffff",
   73941 => x"ffffff",
   73942 => x"ffffff",
   73943 => x"ffffff",
   73944 => x"ffffff",
   73945 => x"ffffff",
   73946 => x"ffffff",
   73947 => x"ffffff",
   73948 => x"ffffff",
   73949 => x"ffffff",
   73950 => x"ffffff",
   73951 => x"ffffff",
   73952 => x"ffffff",
   73953 => x"ffffff",
   73954 => x"ffffff",
   73955 => x"ffffff",
   73956 => x"ffffff",
   73957 => x"ffffff",
   73958 => x"ffffff",
   73959 => x"ffffff",
   73960 => x"ffffff",
   73961 => x"ffffff",
   73962 => x"ffffff",
   73963 => x"ffffff",
   73964 => x"ffffff",
   73965 => x"ffffff",
   73966 => x"ffffff",
   73967 => x"ffffff",
   73968 => x"ffffff",
   73969 => x"ffffff",
   73970 => x"ffffff",
   73971 => x"ffffff",
   73972 => x"ffffff",
   73973 => x"ffffff",
   73974 => x"ffffff",
   73975 => x"ffffff",
   73976 => x"ffffff",
   73977 => x"ffffff",
   73978 => x"ffffff",
   73979 => x"ffffff",
   73980 => x"ffffff",
   73981 => x"ffffff",
   73982 => x"ffffff",
   73983 => x"ffffff",
   73984 => x"ffffff",
   73985 => x"ffffff",
   73986 => x"ffffff",
   73987 => x"ffffff",
   73988 => x"ffffff",
   73989 => x"ffffff",
   73990 => x"ffffff",
   73991 => x"ffffff",
   73992 => x"ffffff",
   73993 => x"ffffff",
   73994 => x"ffffff",
   73995 => x"ffffff",
   73996 => x"ffffff",
   73997 => x"ffffff",
   73998 => x"ffffff",
   73999 => x"ffffff",
   74000 => x"ffffff",
   74001 => x"ffffff",
   74002 => x"ffffff",
   74003 => x"ffffff",
   74004 => x"ffffff",
   74005 => x"ffffff",
   74006 => x"ffffff",
   74007 => x"ffffff",
   74008 => x"ffffff",
   74009 => x"ffffff",
   74010 => x"ffffff",
   74011 => x"ffffff",
   74012 => x"ffffff",
   74013 => x"ffffff",
   74014 => x"ffffff",
   74015 => x"ffffff",
   74016 => x"ffffff",
   74017 => x"ffffff",
   74018 => x"ffffff",
   74019 => x"ffffff",
   74020 => x"ffffff",
   74021 => x"ffffff",
   74022 => x"ffffff",
   74023 => x"ffffff",
   74024 => x"ffffff",
   74025 => x"ffffff",
   74026 => x"ffffff",
   74027 => x"ffffff",
   74028 => x"ffffff",
   74029 => x"ffffff",
   74030 => x"ffffff",
   74031 => x"ffffff",
   74032 => x"ffffff",
   74033 => x"ffffff",
   74034 => x"ffffff",
   74035 => x"ffffff",
   74036 => x"ffffff",
   74037 => x"ffffff",
   74038 => x"ffffff",
   74039 => x"ffffff",
   74040 => x"ffffff",
   74041 => x"ffffff",
   74042 => x"ffffff",
   74043 => x"ffffff",
   74044 => x"ffffff",
   74045 => x"ffffff",
   74046 => x"ffffff",
   74047 => x"ffffff",
   74048 => x"ffffff",
   74049 => x"ffffff",
   74050 => x"ffffff",
   74051 => x"ffffff",
   74052 => x"ffffff",
   74053 => x"ffffff",
   74054 => x"ffffff",
   74055 => x"ffffff",
   74056 => x"ffffff",
   74057 => x"ffffff",
   74058 => x"ffffff",
   74059 => x"ffffff",
   74060 => x"ffffff",
   74061 => x"ffffff",
   74062 => x"ffffff",
   74063 => x"ffffff",
   74064 => x"ffffff",
   74065 => x"ffffff",
   74066 => x"ffffff",
   74067 => x"ffffff",
   74068 => x"ffffff",
   74069 => x"ffffff",
   74070 => x"ffffff",
   74071 => x"ffffff",
   74072 => x"ffffff",
   74073 => x"ffffff",
   74074 => x"ffffff",
   74075 => x"ffffff",
   74076 => x"ffffff",
   74077 => x"ffffff",
   74078 => x"ffffff",
   74079 => x"ffffff",
   74080 => x"ffffff",
   74081 => x"ffffff",
   74082 => x"ffffff",
   74083 => x"ffffff",
   74084 => x"ffffff",
   74085 => x"ffffff",
   74086 => x"ffffff",
   74087 => x"ffffff",
   74088 => x"ffffff",
   74089 => x"ffffff",
   74090 => x"ffffff",
   74091 => x"ffffff",
   74092 => x"ffffff",
   74093 => x"ffffff",
   74094 => x"ffffff",
   74095 => x"ffffff",
   74096 => x"ffffff",
   74097 => x"ffffff",
   74098 => x"ffffff",
   74099 => x"ffffff",
   74100 => x"ffffff",
   74101 => x"ffffff",
   74102 => x"ffffff",
   74103 => x"ffffff",
   74104 => x"ffffff",
   74105 => x"ffffff",
   74106 => x"ffffff",
   74107 => x"ffffff",
   74108 => x"ffffff",
   74109 => x"ffffff",
   74110 => x"ffffff",
   74111 => x"ffffff",
   74112 => x"ffffff",
   74113 => x"ffffff",
   74114 => x"ffffff",
   74115 => x"ffffff",
   74116 => x"ffffff",
   74117 => x"ffffff",
   74118 => x"ffffff",
   74119 => x"ffffff",
   74120 => x"ffffff",
   74121 => x"ffffff",
   74122 => x"ffffff",
   74123 => x"ffffff",
   74124 => x"ffffff",
   74125 => x"ffffff",
   74126 => x"ffffff",
   74127 => x"ffffff",
   74128 => x"ffffff",
   74129 => x"ffffff",
   74130 => x"ffffff",
   74131 => x"ffffff",
   74132 => x"ffffff",
   74133 => x"ffffff",
   74134 => x"ffffff",
   74135 => x"ffffff",
   74136 => x"ffffff",
   74137 => x"ffffff",
   74138 => x"ffffff",
   74139 => x"ffffff",
   74140 => x"ffffff",
   74141 => x"ffffff",
   74142 => x"ffffff",
   74143 => x"ffffff",
   74144 => x"ffffff",
   74145 => x"ffffff",
   74146 => x"ffffff",
   74147 => x"ffffff",
   74148 => x"ffffff",
   74149 => x"ffffff",
   74150 => x"ffffff",
   74151 => x"ffffff",
   74152 => x"ffffff",
   74153 => x"ffffff",
   74154 => x"ffffff",
   74155 => x"ffffff",
   74156 => x"ffffff",
   74157 => x"ffffff",
   74158 => x"ffffff",
   74159 => x"ffffff",
   74160 => x"ffffff",
   74161 => x"ffffff",
   74162 => x"ffffff",
   74163 => x"ffffff",
   74164 => x"ffffff",
   74165 => x"ffffff",
   74166 => x"ffffff",
   74167 => x"ffffff",
   74168 => x"ffffff",
   74169 => x"ffffff",
   74170 => x"ffffff",
   74171 => x"ffffff",
   74172 => x"ffffff",
   74173 => x"ffffff",
   74174 => x"ffffff",
   74175 => x"ffffff",
   74176 => x"ffffff",
   74177 => x"ffffff",
   74178 => x"ffffff",
   74179 => x"ffffff",
   74180 => x"ffffff",
   74181 => x"ffffff",
   74182 => x"ffffff",
   74183 => x"ffffff",
   74184 => x"ffffff",
   74185 => x"ffffff",
   74186 => x"ffffff",
   74187 => x"ffffff",
   74188 => x"ffffff",
   74189 => x"ffffff",
   74190 => x"ffffff",
   74191 => x"ffffff",
   74192 => x"ffffff",
   74193 => x"ffffff",
   74194 => x"ffffff",
   74195 => x"ffffff",
   74196 => x"ffffff",
   74197 => x"ffffff",
   74198 => x"ffffff",
   74199 => x"ffffff",
   74200 => x"ffffff",
   74201 => x"ffffff",
   74202 => x"ffffff",
   74203 => x"ffffff",
   74204 => x"ffffff",
   74205 => x"ffffff",
   74206 => x"ffffff",
   74207 => x"ffffff",
   74208 => x"ffffff",
   74209 => x"ffffff",
   74210 => x"ffffff",
   74211 => x"ffffff",
   74212 => x"ffffff",
   74213 => x"ffffff",
   74214 => x"ffffff",
   74215 => x"ffffff",
   74216 => x"ffffff",
   74217 => x"ffffff",
   74218 => x"ffffff",
   74219 => x"ffffff",
   74220 => x"ffffff",
   74221 => x"ffffff",
   74222 => x"ffffff",
   74223 => x"ffffff",
   74224 => x"ffffff",
   74225 => x"ffffff",
   74226 => x"ffffff",
   74227 => x"ffffff",
   74228 => x"ffffff",
   74229 => x"ffffff",
   74230 => x"ffffff",
   74231 => x"ffffff",
   74232 => x"ffffff",
   74233 => x"ffffff",
   74234 => x"ffffff",
   74235 => x"ffffff",
   74236 => x"ffffff",
   74237 => x"ffffff",
   74238 => x"ffffff",
   74239 => x"ffffff",
   74240 => x"ffffff",
   74241 => x"ffffff",
   74242 => x"ffffff",
   74243 => x"ffffff",
   74244 => x"ffffff",
   74245 => x"ffffff",
   74246 => x"ffffff",
   74247 => x"ffffff",
   74248 => x"ffffff",
   74249 => x"ffffff",
   74250 => x"ffffff",
   74251 => x"ffffff",
   74252 => x"ffffff",
   74253 => x"ffffff",
   74254 => x"ffffff",
   74255 => x"ffffff",
   74256 => x"ffffff",
   74257 => x"ffffff",
   74258 => x"ffffff",
   74259 => x"ffffff",
   74260 => x"ffffff",
   74261 => x"ffffff",
   74262 => x"ffffff",
   74263 => x"ffffff",
   74264 => x"ffffff",
   74265 => x"ffffff",
   74266 => x"ffffff",
   74267 => x"ffffff",
   74268 => x"ffffff",
   74269 => x"ffffff",
   74270 => x"ffffff",
   74271 => x"ffffff",
   74272 => x"ffffff",
   74273 => x"ffffff",
   74274 => x"ffffff",
   74275 => x"ffffff",
   74276 => x"ffffff",
   74277 => x"ffffff",
   74278 => x"ffffff",
   74279 => x"ffffff",
   74280 => x"ffffff",
   74281 => x"ffffff",
   74282 => x"ffffff",
   74283 => x"ffffff",
   74284 => x"ffffff",
   74285 => x"ffffff",
   74286 => x"ffffff",
   74287 => x"ffffff",
   74288 => x"ffffff",
   74289 => x"ffffff",
   74290 => x"ffffff",
   74291 => x"ffffff",
   74292 => x"ffffff",
   74293 => x"ffffff",
   74294 => x"ffffff",
   74295 => x"ffffff",
   74296 => x"ffffff",
   74297 => x"ffffff",
   74298 => x"ffffff",
   74299 => x"ffffff",
   74300 => x"ffffff",
   74301 => x"ffffff",
   74302 => x"ffffff",
   74303 => x"ffffff",
   74304 => x"ffffff",
   74305 => x"ffffff",
   74306 => x"ffffff",
   74307 => x"ffffff",
   74308 => x"ffffff",
   74309 => x"ffffff",
   74310 => x"ffffff",
   74311 => x"ffffff",
   74312 => x"ffffff",
   74313 => x"ffffff",
   74314 => x"ffffff",
   74315 => x"ffffff",
   74316 => x"ffffff",
   74317 => x"ffffff",
   74318 => x"ffffff",
   74319 => x"ffffff",
   74320 => x"ffffff",
   74321 => x"ffffff",
   74322 => x"ffffff",
   74323 => x"ffffff",
   74324 => x"ffffff",
   74325 => x"ffffff",
   74326 => x"ffffff",
   74327 => x"ffffff",
   74328 => x"ffffff",
   74329 => x"ffffff",
   74330 => x"ffffff",
   74331 => x"ffffff",
   74332 => x"ffffff",
   74333 => x"ffffff",
   74334 => x"ffffff",
   74335 => x"ffffff",
   74336 => x"ffffff",
   74337 => x"ffffff",
   74338 => x"ffffff",
   74339 => x"ffffff",
   74340 => x"ffffff",
   74341 => x"ffffff",
   74342 => x"ffffff",
   74343 => x"ffffff",
   74344 => x"ffffff",
   74345 => x"ffffff",
   74346 => x"ffffff",
   74347 => x"ffffff",
   74348 => x"ffffff",
   74349 => x"ffffff",
   74350 => x"ffffff",
   74351 => x"ffffff",
   74352 => x"ffffff",
   74353 => x"ffffff",
   74354 => x"ffffff",
   74355 => x"ffffff",
   74356 => x"ffffff",
   74357 => x"ffffff",
   74358 => x"ffffff",
   74359 => x"ffffff",
   74360 => x"ffffff",
   74361 => x"ffffff",
   74362 => x"ffffff",
   74363 => x"ffffff",
   74364 => x"ffffff",
   74365 => x"ffffff",
   74366 => x"ffffff",
   74367 => x"ffffff",
   74368 => x"ffffff",
   74369 => x"ffffff",
   74370 => x"ffffff",
   74371 => x"ffffff",
   74372 => x"ffffff",
   74373 => x"ffffff",
   74374 => x"ffffff",
   74375 => x"ffffff",
   74376 => x"ffffff",
   74377 => x"ffffff",
   74378 => x"ffffff",
   74379 => x"ffffff",
   74380 => x"ffffff",
   74381 => x"ffffff",
   74382 => x"ffffff",
   74383 => x"ffffff",
   74384 => x"ffffff",
   74385 => x"ffffff",
   74386 => x"ffffff",
   74387 => x"ffffff",
   74388 => x"ffffff",
   74389 => x"ffffff",
   74390 => x"ffffff",
   74391 => x"ffffff",
   74392 => x"ffffff",
   74393 => x"ffffff",
   74394 => x"ffffff",
   74395 => x"ffffff",
   74396 => x"ffffff",
   74397 => x"ffffff",
   74398 => x"ffffff",
   74399 => x"ffffff",
   74400 => x"ffffff",
   74401 => x"ffffff",
   74402 => x"ffffff",
   74403 => x"ffffff",
   74404 => x"ffffff",
   74405 => x"ffffff",
   74406 => x"ffffff",
   74407 => x"ffffff",
   74408 => x"ffffff",
   74409 => x"ffffff",
   74410 => x"ffffff",
   74411 => x"ffffff",
   74412 => x"ffffff",
   74413 => x"ffffff",
   74414 => x"ffffff",
   74415 => x"ffffff",
   74416 => x"ffffff",
   74417 => x"ffffff",
   74418 => x"ffffff",
   74419 => x"ffffff",
   74420 => x"ffffff",
   74421 => x"ffffff",
   74422 => x"ffffff",
   74423 => x"ffffff",
   74424 => x"ffffff",
   74425 => x"ffffff",
   74426 => x"ffffff",
   74427 => x"ffffff",
   74428 => x"ffffff",
   74429 => x"ffffff",
   74430 => x"ffffff",
   74431 => x"ffffff",
   74432 => x"ffffff",
   74433 => x"ffffff",
   74434 => x"ffffff",
   74435 => x"ffffff",
   74436 => x"ffffff",
   74437 => x"ffffff",
   74438 => x"ffffff",
   74439 => x"ffffff",
   74440 => x"ffffff",
   74441 => x"ffffff",
   74442 => x"ffffff",
   74443 => x"ffffff",
   74444 => x"ffffff",
   74445 => x"ffffff",
   74446 => x"ffffff",
   74447 => x"ffffff",
   74448 => x"ffffff",
   74449 => x"ffffff",
   74450 => x"ffffff",
   74451 => x"ffffff",
   74452 => x"ffffff",
   74453 => x"ffffff",
   74454 => x"ffffff",
   74455 => x"ffffff",
   74456 => x"ffffff",
   74457 => x"ffffff",
   74458 => x"ffffff",
   74459 => x"ffffff",
   74460 => x"ffffff",
   74461 => x"ffffff",
   74462 => x"ffffff",
   74463 => x"ffffff",
   74464 => x"ffffff",
   74465 => x"ffffff",
   74466 => x"ffffff",
   74467 => x"ffffff",
   74468 => x"ffffff",
   74469 => x"ffffff",
   74470 => x"ffffff",
   74471 => x"ffffff",
   74472 => x"ffffff",
   74473 => x"ffffff",
   74474 => x"ffffff",
   74475 => x"ffffff",
   74476 => x"ffffff",
   74477 => x"ffffff",
   74478 => x"ffffff",
   74479 => x"ffffff",
   74480 => x"ffffff",
   74481 => x"ffffff",
   74482 => x"ffffff",
   74483 => x"ffffff",
   74484 => x"ffffff",
   74485 => x"ffffff",
   74486 => x"ffffff",
   74487 => x"ffffff",
   74488 => x"ffffff",
   74489 => x"ffffff",
   74490 => x"ffffff",
   74491 => x"ffffff",
   74492 => x"ffffff",
   74493 => x"ffffff",
   74494 => x"ffffff",
   74495 => x"ffffff",
   74496 => x"ffffff",
   74497 => x"ffffff",
   74498 => x"ffffff",
   74499 => x"ffffff",
   74500 => x"ffffff",
   74501 => x"ffffff",
   74502 => x"ffffff",
   74503 => x"ffffff",
   74504 => x"ffffff",
   74505 => x"ffffff",
   74506 => x"ffffff",
   74507 => x"ffffff",
   74508 => x"ffffff",
   74509 => x"ffffff",
   74510 => x"ffffff",
   74511 => x"ffffff",
   74512 => x"ffffff",
   74513 => x"ffffff",
   74514 => x"ffffff",
   74515 => x"ffffff",
   74516 => x"ffffff",
   74517 => x"ffffff",
   74518 => x"ffffff",
   74519 => x"ffffff",
   74520 => x"ffffff",
   74521 => x"ffffff",
   74522 => x"ffffff",
   74523 => x"ffffff",
   74524 => x"ffffff",
   74525 => x"ffffff",
   74526 => x"ffffff",
   74527 => x"ffffff",
   74528 => x"ffffff",
   74529 => x"ffffff",
   74530 => x"ffffff",
   74531 => x"ffffff",
   74532 => x"ffffff",
   74533 => x"ffffff",
   74534 => x"ffffff",
   74535 => x"ffffff",
   74536 => x"ffffff",
   74537 => x"ffffff",
   74538 => x"ffffff",
   74539 => x"ffffff",
   74540 => x"ffffff",
   74541 => x"ffffff",
   74542 => x"ffffff",
   74543 => x"ffffff",
   74544 => x"ffffff",
   74545 => x"ffffff",
   74546 => x"ffffff",
   74547 => x"ffffff",
   74548 => x"ffffff",
   74549 => x"ffffff",
   74550 => x"ffffff",
   74551 => x"ffffff",
   74552 => x"ffffff",
   74553 => x"ffffff",
   74554 => x"ffffff",
   74555 => x"ffffff",
   74556 => x"ffffff",
   74557 => x"ffffff",
   74558 => x"ffffff",
   74559 => x"ffffff",
   74560 => x"ffffff",
   74561 => x"ffffff",
   74562 => x"ffffff",
   74563 => x"ffffff",
   74564 => x"ffffff",
   74565 => x"ffffff",
   74566 => x"ffffff",
   74567 => x"ffffff",
   74568 => x"ffffff",
   74569 => x"ffffff",
   74570 => x"ffffff",
   74571 => x"ffffff",
   74572 => x"ffffff",
   74573 => x"ffffff",
   74574 => x"ffffff",
   74575 => x"ffffff",
   74576 => x"ffffff",
   74577 => x"ffffff",
   74578 => x"ffffff",
   74579 => x"ffffff",
   74580 => x"ffffff",
   74581 => x"ffffff",
   74582 => x"ffffff",
   74583 => x"ffffff",
   74584 => x"ffffff",
   74585 => x"ffffff",
   74586 => x"ffffff",
   74587 => x"ffffff",
   74588 => x"ffffff",
   74589 => x"ffffff",
   74590 => x"ffffff",
   74591 => x"ffffff",
   74592 => x"ffffff",
   74593 => x"ffffff",
   74594 => x"ffffff",
   74595 => x"ffffff",
   74596 => x"ffffff",
   74597 => x"ffffff",
   74598 => x"ffffff",
   74599 => x"ffffff",
   74600 => x"ffffff",
   74601 => x"ffffff",
   74602 => x"ffffff",
   74603 => x"ffffff",
   74604 => x"ffffff",
   74605 => x"ffffff",
   74606 => x"ffffff",
   74607 => x"ffffff",
   74608 => x"ffffff",
   74609 => x"ffffff",
   74610 => x"ffffff",
   74611 => x"ffffff",
   74612 => x"ffffff",
   74613 => x"ffffff",
   74614 => x"ffffff",
   74615 => x"ffffff",
   74616 => x"ffffff",
   74617 => x"ffffff",
   74618 => x"ffffff",
   74619 => x"ffffff",
   74620 => x"ffffff",
   74621 => x"ffffff",
   74622 => x"ffffff",
   74623 => x"ffffff",
   74624 => x"ffffff",
   74625 => x"ffffff",
   74626 => x"ffffff",
   74627 => x"ffffff",
   74628 => x"ffffff",
   74629 => x"ffffff",
   74630 => x"ffffff",
   74631 => x"ffffff",
   74632 => x"ffffff",
   74633 => x"ffffff",
   74634 => x"ffffff",
   74635 => x"ffffff",
   74636 => x"ffffff",
   74637 => x"ffffff",
   74638 => x"ffffff",
   74639 => x"ffffff",
   74640 => x"ffffff",
   74641 => x"ffffff",
   74642 => x"ffffff",
   74643 => x"ffffff",
   74644 => x"ffffff",
   74645 => x"ffffff",
   74646 => x"ffffff",
   74647 => x"ffffff",
   74648 => x"ffffff",
   74649 => x"ffffff",
   74650 => x"ffffff",
   74651 => x"ffffff",
   74652 => x"ffffff",
   74653 => x"ffffff",
   74654 => x"ffffff",
   74655 => x"ffffff",
   74656 => x"ffffff",
   74657 => x"ffffff",
   74658 => x"ffffff",
   74659 => x"ffffff",
   74660 => x"ffffff",
   74661 => x"ffffff",
   74662 => x"ffffff",
   74663 => x"ffffff",
   74664 => x"ffffff",
   74665 => x"ffffff",
   74666 => x"ffffff",
   74667 => x"ffffff",
   74668 => x"ffffff",
   74669 => x"ffffff",
   74670 => x"ffffff",
   74671 => x"ffffff",
   74672 => x"ffffff",
   74673 => x"ffffff",
   74674 => x"ffffff",
   74675 => x"ffffff",
   74676 => x"ffffff",
   74677 => x"ffffff",
   74678 => x"ffffff",
   74679 => x"ffffff",
   74680 => x"ffffff",
   74681 => x"ffffff",
   74682 => x"ffffff",
   74683 => x"ffffff",
   74684 => x"ffffff",
   74685 => x"ffffff",
   74686 => x"ffffff",
   74687 => x"ffffff",
   74688 => x"ffffff",
   74689 => x"ffffff",
   74690 => x"ffffff",
   74691 => x"ffffff",
   74692 => x"ffffff",
   74693 => x"ffffff",
   74694 => x"ffffff",
   74695 => x"ffffff",
   74696 => x"ffffff",
   74697 => x"ffffff",
   74698 => x"ffffff",
   74699 => x"ffffff",
   74700 => x"ffffff",
   74701 => x"ffffff",
   74702 => x"ffffff",
   74703 => x"ffffff",
   74704 => x"ffffff",
   74705 => x"ffffff",
   74706 => x"ffffff",
   74707 => x"ffffff",
   74708 => x"ffffff",
   74709 => x"ffffff",
   74710 => x"ffffff",
   74711 => x"ffffff",
   74712 => x"ffffff",
   74713 => x"ffffff",
   74714 => x"ffffff",
   74715 => x"ffffff",
   74716 => x"ffffff",
   74717 => x"ffffff",
   74718 => x"ffffff",
   74719 => x"ffffff",
   74720 => x"ffffff",
   74721 => x"ffffff",
   74722 => x"ffffff",
   74723 => x"ffffff",
   74724 => x"ffffff",
   74725 => x"ffffff",
   74726 => x"ffffff",
   74727 => x"ffffff",
   74728 => x"ffffff",
   74729 => x"ffffff",
   74730 => x"ffffff",
   74731 => x"ffffff",
   74732 => x"ffffff",
   74733 => x"ffffff",
   74734 => x"ffffff",
   74735 => x"ffffff",
   74736 => x"ffffff",
   74737 => x"ffffff",
   74738 => x"ffffff",
   74739 => x"ffffff",
   74740 => x"ffffff",
   74741 => x"ffffff",
   74742 => x"ffffff",
   74743 => x"ffffff",
   74744 => x"ffffff",
   74745 => x"ffffff",
   74746 => x"ffffff",
   74747 => x"ffffff",
   74748 => x"ffffff",
   74749 => x"ffffff",
   74750 => x"ffffff",
   74751 => x"ffffff",
   74752 => x"ffffff",
   74753 => x"ffffff",
   74754 => x"ffffff",
   74755 => x"ffffff",
   74756 => x"ffffff",
   74757 => x"ffffff",
   74758 => x"ffffff",
   74759 => x"ffffff",
   74760 => x"ffffff",
   74761 => x"ffffff",
   74762 => x"ffffff",
   74763 => x"ffffff",
   74764 => x"ffffff",
   74765 => x"ffffff",
   74766 => x"ffffff",
   74767 => x"ffffff",
   74768 => x"ffffff",
   74769 => x"ffffff",
   74770 => x"ffffff",
   74771 => x"ffffff",
   74772 => x"ffffff",
   74773 => x"ffffff",
   74774 => x"ffffff",
   74775 => x"ffffff",
   74776 => x"ffffff",
   74777 => x"ffffff",
   74778 => x"ffffff",
   74779 => x"ffffff",
   74780 => x"ffffff",
   74781 => x"ffffff",
   74782 => x"ffffff",
   74783 => x"ffffff",
   74784 => x"ffffff",
   74785 => x"ffffff",
   74786 => x"ffffff",
   74787 => x"ffffff",
   74788 => x"ffffff",
   74789 => x"ffffff",
   74790 => x"ffffff",
   74791 => x"ffffff",
   74792 => x"ffffff",
   74793 => x"ffffff",
   74794 => x"ffffff",
   74795 => x"ffffff",
   74796 => x"ffffff",
   74797 => x"ffffff",
   74798 => x"ffffff",
   74799 => x"ffffff",
   74800 => x"ffffff",
   74801 => x"ffffff",
   74802 => x"ffffff",
   74803 => x"ffffff",
   74804 => x"ffffff",
   74805 => x"ffffff",
   74806 => x"ffffff",
   74807 => x"ffffff",
   74808 => x"ffffff",
   74809 => x"ffffff",
   74810 => x"ffffff",
   74811 => x"ffffff",
   74812 => x"ffffff",
   74813 => x"ffffff",
   74814 => x"ffffff",
   74815 => x"ffffff",
   74816 => x"ffffff",
   74817 => x"ffffff",
   74818 => x"ffffff",
   74819 => x"ffffff",
   74820 => x"ffffff",
   74821 => x"ffffff",
   74822 => x"ffffff",
   74823 => x"ffffff",
   74824 => x"ffffff",
   74825 => x"ffffff",
   74826 => x"ffffff",
   74827 => x"ffffff",
   74828 => x"ffffff",
   74829 => x"ffffff",
   74830 => x"ffffff",
   74831 => x"ffffff",
   74832 => x"ffffff",
   74833 => x"ffffff",
   74834 => x"ffffff",
   74835 => x"ffffff",
   74836 => x"ffffff",
   74837 => x"ffffff",
   74838 => x"ffffff",
   74839 => x"ffffff",
   74840 => x"ffffff",
   74841 => x"ffffff",
   74842 => x"ffffff",
   74843 => x"ffffff",
   74844 => x"ffffff",
   74845 => x"ffffff",
   74846 => x"ffffff",
   74847 => x"ffffff",
   74848 => x"ffffff",
   74849 => x"ffffff",
   74850 => x"ffffff",
   74851 => x"ffffff",
   74852 => x"ffffff",
   74853 => x"ffffff",
   74854 => x"ffffff",
   74855 => x"ffffff",
   74856 => x"ffffff",
   74857 => x"ffffff",
   74858 => x"ffffff",
   74859 => x"ffffff",
   74860 => x"ffffff",
   74861 => x"ffffff",
   74862 => x"ffffff",
   74863 => x"ffffff",
   74864 => x"ffffff",
   74865 => x"ffffff",
   74866 => x"ffffff",
   74867 => x"ffffff",
   74868 => x"ffffff",
   74869 => x"ffffff",
   74870 => x"ffffff",
   74871 => x"ffffff",
   74872 => x"ffffff",
   74873 => x"ffffff",
   74874 => x"ffffff",
   74875 => x"ffffff",
   74876 => x"ffffff",
   74877 => x"ffffff",
   74878 => x"ffffff",
   74879 => x"ffffff",
   74880 => x"ffffff",
   74881 => x"ffffff",
   74882 => x"ffffff",
   74883 => x"ffffff",
   74884 => x"ffffff",
   74885 => x"ffffff",
   74886 => x"ffffff",
   74887 => x"ffffff",
   74888 => x"ffffff",
   74889 => x"ffffff",
   74890 => x"ffffff",
   74891 => x"ffffff",
   74892 => x"ffffff",
   74893 => x"ffffff",
   74894 => x"ffffff",
   74895 => x"ffffff",
   74896 => x"ffffff",
   74897 => x"ffffff",
   74898 => x"ffffff",
   74899 => x"ffffff",
   74900 => x"ffffff",
   74901 => x"ffffff",
   74902 => x"ffffff",
   74903 => x"ffffff",
   74904 => x"ffffff",
   74905 => x"ffffff",
   74906 => x"ffffff",
   74907 => x"ffffff",
   74908 => x"ffffff",
   74909 => x"ffffff",
   74910 => x"ffffff",
   74911 => x"ffffff",
   74912 => x"ffffff",
   74913 => x"ffffff",
   74914 => x"ffffff",
   74915 => x"ffffff",
   74916 => x"ffffff",
   74917 => x"ffffff",
   74918 => x"ffffff",
   74919 => x"ffffff",
   74920 => x"ffffff",
   74921 => x"ffffff",
   74922 => x"ffffff",
   74923 => x"ffffff",
   74924 => x"ffffff",
   74925 => x"ffffff",
   74926 => x"ffffff",
   74927 => x"ffffff",
   74928 => x"ffffff",
   74929 => x"ffffff",
   74930 => x"ffffff",
   74931 => x"ffffff",
   74932 => x"ffffff",
   74933 => x"ffffff",
   74934 => x"ffffff",
   74935 => x"ffffff",
   74936 => x"ffffff",
   74937 => x"ffffff",
   74938 => x"ffffff",
   74939 => x"ffffff",
   74940 => x"ffffff",
   74941 => x"ffffff",
   74942 => x"ffffff",
   74943 => x"ffffff",
   74944 => x"ffffff",
   74945 => x"ffffff",
   74946 => x"ffffff",
   74947 => x"ffffff",
   74948 => x"ffffff",
   74949 => x"ffffff",
   74950 => x"ffffff",
   74951 => x"ffffff",
   74952 => x"ffffff",
   74953 => x"ffffff",
   74954 => x"ffffff",
   74955 => x"ffffff",
   74956 => x"ffffff",
   74957 => x"ffffff",
   74958 => x"ffffff",
   74959 => x"ffffff",
   74960 => x"ffffff",
   74961 => x"ffffff",
   74962 => x"ffffff",
   74963 => x"ffffff",
   74964 => x"ffffff",
   74965 => x"ffffff",
   74966 => x"ffffff",
   74967 => x"ffffff",
   74968 => x"ffffff",
   74969 => x"ffffff",
   74970 => x"ffffff",
   74971 => x"ffffff",
   74972 => x"ffffff",
   74973 => x"ffffff",
   74974 => x"ffffff",
   74975 => x"ffffff",
   74976 => x"ffffff",
   74977 => x"ffffff",
   74978 => x"ffffff",
   74979 => x"ffffff",
   74980 => x"ffffff",
   74981 => x"ffffff",
   74982 => x"ffffff",
   74983 => x"ffffff",
   74984 => x"ffffff",
   74985 => x"ffffff",
   74986 => x"ffffff",
   74987 => x"ffffff",
   74988 => x"ffffff",
   74989 => x"ffffff",
   74990 => x"ffffff",
   74991 => x"ffffff",
   74992 => x"ffffff",
   74993 => x"ffffff",
   74994 => x"ffffff",
   74995 => x"ffffff",
   74996 => x"ffffff",
   74997 => x"ffffff",
   74998 => x"ffffff",
   74999 => x"ffffff",
   75000 => x"ffffff",
   75001 => x"ffffff",
   75002 => x"ffffff",
   75003 => x"ffffff",
   75004 => x"ffffff",
   75005 => x"ffffff",
   75006 => x"ffffff",
   75007 => x"ffffff",
   75008 => x"ffffff",
   75009 => x"ffffff",
   75010 => x"ffffff",
   75011 => x"ffffff",
   75012 => x"ffffff",
   75013 => x"ffffff",
   75014 => x"ffffff",
   75015 => x"ffffff",
   75016 => x"ffffff",
   75017 => x"ffffff",
   75018 => x"ffffff",
   75019 => x"ffffff",
   75020 => x"ffffff",
   75021 => x"ffffff",
   75022 => x"ffffff",
   75023 => x"ffffff",
   75024 => x"ffffff",
   75025 => x"ffffff",
   75026 => x"ffffff",
   75027 => x"ffffff",
   75028 => x"ffffff",
   75029 => x"ffffff",
   75030 => x"ffffff",
   75031 => x"ffffff",
   75032 => x"ffffff",
   75033 => x"ffffff",
   75034 => x"ffffff",
   75035 => x"ffffff",
   75036 => x"ffffff",
   75037 => x"ffffff",
   75038 => x"ffffff",
   75039 => x"ffffff",
   75040 => x"ffffff",
   75041 => x"ffffff",
   75042 => x"ffffff",
   75043 => x"ffffff",
   75044 => x"ffffff",
   75045 => x"ffffff",
   75046 => x"ffffff",
   75047 => x"ffffff",
   75048 => x"ffffff",
   75049 => x"ffffff",
   75050 => x"ffffff",
   75051 => x"ffffff",
   75052 => x"ffffff",
   75053 => x"ffffff",
   75054 => x"ffffff",
   75055 => x"ffffff",
   75056 => x"ffffff",
   75057 => x"ffffff",
   75058 => x"ffffff",
   75059 => x"ffffff",
   75060 => x"ffffff",
   75061 => x"ffffff",
   75062 => x"ffffff",
   75063 => x"ffffff",
   75064 => x"ffffff",
   75065 => x"ffffff",
   75066 => x"ffffff",
   75067 => x"ffffff",
   75068 => x"ffffff",
   75069 => x"ffffff",
   75070 => x"ffffff",
   75071 => x"ffffff",
   75072 => x"ffffff",
   75073 => x"ffffff",
   75074 => x"ffffff",
   75075 => x"ffffff",
   75076 => x"ffffff",
   75077 => x"ffffff",
   75078 => x"ffffff",
   75079 => x"ffffff",
   75080 => x"ffffff",
   75081 => x"ffffff",
   75082 => x"ffffff",
   75083 => x"ffffff",
   75084 => x"ffffff",
   75085 => x"ffffff",
   75086 => x"ffffff",
   75087 => x"ffffff",
   75088 => x"ffffff",
   75089 => x"ffffff",
   75090 => x"ffffff",
   75091 => x"ffffff",
   75092 => x"ffffff",
   75093 => x"ffffff",
   75094 => x"ffffff",
   75095 => x"ffffff",
   75096 => x"ffffff",
   75097 => x"ffffff",
   75098 => x"ffffff",
   75099 => x"ffffff",
   75100 => x"ffffff",
   75101 => x"ffffff",
   75102 => x"ffffff",
   75103 => x"ffffff",
   75104 => x"ffffff",
   75105 => x"ffffff",
   75106 => x"ffffff",
   75107 => x"ffffff",
   75108 => x"ffffff",
   75109 => x"ffffff",
   75110 => x"ffffff",
   75111 => x"ffffff",
   75112 => x"ffffff",
   75113 => x"ffffff",
   75114 => x"ffffff",
   75115 => x"ffffff",
   75116 => x"ffffff",
   75117 => x"ffffff",
   75118 => x"ffffff",
   75119 => x"ffffff",
   75120 => x"ffffff",
   75121 => x"ffffff",
   75122 => x"ffffff",
   75123 => x"ffffff",
   75124 => x"ffffff",
   75125 => x"ffffff",
   75126 => x"ffffff",
   75127 => x"ffffff",
   75128 => x"ffffff",
   75129 => x"ffffff",
   75130 => x"ffffff",
   75131 => x"ffffff",
   75132 => x"ffffff",
   75133 => x"ffffff",
   75134 => x"ffffff",
   75135 => x"ffffff",
   75136 => x"ffffff",
   75137 => x"ffffff",
   75138 => x"ffffff",
   75139 => x"ffffff",
   75140 => x"ffffff",
   75141 => x"ffffff",
   75142 => x"ffffff",
   75143 => x"ffffff",
   75144 => x"ffffff",
   75145 => x"ffffff",
   75146 => x"ffffff",
   75147 => x"ffffff",
   75148 => x"ffffff",
   75149 => x"ffffff",
   75150 => x"ffffff",
   75151 => x"ffffff",
   75152 => x"ffffff",
   75153 => x"ffffff",
   75154 => x"ffffff",
   75155 => x"ffffff",
   75156 => x"ffffff",
   75157 => x"ffffff",
   75158 => x"ffffff",
   75159 => x"ffffff",
   75160 => x"ffffff",
   75161 => x"ffffff",
   75162 => x"ffffff",
   75163 => x"ffffff",
   75164 => x"ffffff",
   75165 => x"ffffff",
   75166 => x"ffffff",
   75167 => x"ffffff",
   75168 => x"ffffff",
   75169 => x"ffffff",
   75170 => x"ffffff",
   75171 => x"ffffff",
   75172 => x"ffffff",
   75173 => x"ffffff",
   75174 => x"ffffff",
   75175 => x"ffffff",
   75176 => x"ffffff",
   75177 => x"ffffff",
   75178 => x"ffffff",
   75179 => x"ffffff",
   75180 => x"ffffff",
   75181 => x"ffffff",
   75182 => x"ffffff",
   75183 => x"ffffff",
   75184 => x"ffffff",
   75185 => x"ffffff",
   75186 => x"ffffff",
   75187 => x"ffffff",
   75188 => x"ffffff",
   75189 => x"ffffff",
   75190 => x"ffffff",
   75191 => x"ffffff",
   75192 => x"ffffff",
   75193 => x"ffffff",
   75194 => x"ffffff",
   75195 => x"ffffff",
   75196 => x"ffffff",
   75197 => x"ffffff",
   75198 => x"ffffff",
   75199 => x"ffffff",
   75200 => x"ffffff",
   75201 => x"ffffff",
   75202 => x"ffffff",
   75203 => x"ffffff",
   75204 => x"ffffff",
   75205 => x"ffffff",
   75206 => x"ffffff",
   75207 => x"ffffff",
   75208 => x"ffffff",
   75209 => x"ffffff",
   75210 => x"ffffff",
   75211 => x"ffffff",
   75212 => x"ffffff",
   75213 => x"ffffff",
   75214 => x"ffffff",
   75215 => x"ffffff",
   75216 => x"ffffff",
   75217 => x"ffffff",
   75218 => x"ffffff",
   75219 => x"ffffff",
   75220 => x"ffffff",
   75221 => x"ffffff",
   75222 => x"ffffff",
   75223 => x"ffffff",
   75224 => x"ffffff",
   75225 => x"ffffff",
   75226 => x"ffffff",
   75227 => x"ffffff",
   75228 => x"ffffff",
   75229 => x"ffffff",
   75230 => x"ffffff",
   75231 => x"ffffff",
   75232 => x"ffffff",
   75233 => x"ffffff",
   75234 => x"ffffff",
   75235 => x"ffffff",
   75236 => x"ffffff",
   75237 => x"ffffff",
   75238 => x"ffffff",
   75239 => x"ffffff",
   75240 => x"ffffff",
   75241 => x"ffffff",
   75242 => x"ffffff",
   75243 => x"ffffff",
   75244 => x"ffffff",
   75245 => x"ffffff",
   75246 => x"ffffff",
   75247 => x"ffffff",
   75248 => x"ffffff",
   75249 => x"ffffff",
   75250 => x"ffffff",
   75251 => x"ffffff",
   75252 => x"ffffff",
   75253 => x"ffffff",
   75254 => x"ffffff",
   75255 => x"ffffff",
   75256 => x"ffffff",
   75257 => x"ffffff",
   75258 => x"ffffff",
   75259 => x"ffffff",
   75260 => x"ffffff",
   75261 => x"ffffff",
   75262 => x"ffffff",
   75263 => x"ffffff",
   75264 => x"ffffff",
   75265 => x"ffffff",
   75266 => x"ffffff",
   75267 => x"ffffff",
   75268 => x"ffffff",
   75269 => x"ffffff",
   75270 => x"ffffff",
   75271 => x"ffffff",
   75272 => x"ffffff",
   75273 => x"ffffff",
   75274 => x"ffffff",
   75275 => x"ffffff",
   75276 => x"ffffff",
   75277 => x"ffffff",
   75278 => x"ffffff",
   75279 => x"ffffff",
   75280 => x"ffffff",
   75281 => x"ffffff",
   75282 => x"ffffff",
   75283 => x"ffffff",
   75284 => x"ffffff",
   75285 => x"ffffff",
   75286 => x"ffffff",
   75287 => x"ffffff",
   75288 => x"ffffff",
   75289 => x"ffffff",
   75290 => x"ffffff",
   75291 => x"ffffff",
   75292 => x"ffffff",
   75293 => x"ffffff",
   75294 => x"ffffff",
   75295 => x"ffffff",
   75296 => x"ffffff",
   75297 => x"ffffff",
   75298 => x"ffffff",
   75299 => x"ffffff",
   75300 => x"ffffff",
   75301 => x"ffffff",
   75302 => x"ffffff",
   75303 => x"ffffff",
   75304 => x"ffffff",
   75305 => x"ffffff",
   75306 => x"ffffff",
   75307 => x"ffffff",
   75308 => x"ffffff",
   75309 => x"ffffff",
   75310 => x"ffffff",
   75311 => x"ffffff",
   75312 => x"ffffff",
   75313 => x"ffffff",
   75314 => x"ffffff",
   75315 => x"ffffff",
   75316 => x"ffffff",
   75317 => x"ffffff",
   75318 => x"ffffff",
   75319 => x"ffffff",
   75320 => x"ffffff",
   75321 => x"ffffff",
   75322 => x"ffffff",
   75323 => x"ffffff",
   75324 => x"ffffff",
   75325 => x"ffffff",
   75326 => x"ffffff",
   75327 => x"ffffff",
   75328 => x"ffffff",
   75329 => x"ffffff",
   75330 => x"ffffff",
   75331 => x"ffffff",
   75332 => x"ffffff",
   75333 => x"ffffff",
   75334 => x"ffffff",
   75335 => x"ffffff",
   75336 => x"ffffff",
   75337 => x"ffffff",
   75338 => x"ffffff",
   75339 => x"ffffff",
   75340 => x"ffffff",
   75341 => x"ffffff",
   75342 => x"ffffff",
   75343 => x"ffffff",
   75344 => x"ffffff",
   75345 => x"ffffff",
   75346 => x"ffffff",
   75347 => x"ffffff",
   75348 => x"ffffff",
   75349 => x"ffffff",
   75350 => x"ffffff",
   75351 => x"ffffff",
   75352 => x"ffffff",
   75353 => x"ffffff",
   75354 => x"ffffff",
   75355 => x"ffffff",
   75356 => x"ffffff",
   75357 => x"ffffff",
   75358 => x"ffffff",
   75359 => x"ffffff",
   75360 => x"ffffff",
   75361 => x"ffffff",
   75362 => x"ffffff",
   75363 => x"ffffff",
   75364 => x"ffffff",
   75365 => x"ffffff",
   75366 => x"ffffff",
   75367 => x"ffffff",
   75368 => x"ffffff",
   75369 => x"ffffff",
   75370 => x"ffffff",
   75371 => x"ffffff",
   75372 => x"ffffff",
   75373 => x"ffffff",
   75374 => x"ffffff",
   75375 => x"ffffff",
   75376 => x"ffffff",
   75377 => x"ffffff",
   75378 => x"ffffff",
   75379 => x"ffffff",
   75380 => x"ffffff",
   75381 => x"ffffff",
   75382 => x"ffffff",
   75383 => x"ffffff",
   75384 => x"ffffff",
   75385 => x"ffffff",
   75386 => x"ffffff",
   75387 => x"ffffff",
   75388 => x"ffffff",
   75389 => x"ffffff",
   75390 => x"ffffff",
   75391 => x"ffffff",
   75392 => x"ffffff",
   75393 => x"ffffff",
   75394 => x"ffffff",
   75395 => x"ffffff",
   75396 => x"ffffff",
   75397 => x"ffffff",
   75398 => x"ffffff",
   75399 => x"ffffff",
   75400 => x"ffffff",
   75401 => x"ffffff",
   75402 => x"ffffff",
   75403 => x"ffffff",
   75404 => x"ffffff",
   75405 => x"ffffff",
   75406 => x"ffffff",
   75407 => x"ffffff",
   75408 => x"ffffff",
   75409 => x"ffffff",
   75410 => x"ffffff",
   75411 => x"ffffff",
   75412 => x"ffffff",
   75413 => x"ffffff",
   75414 => x"ffffff",
   75415 => x"ffffff",
   75416 => x"ffffff",
   75417 => x"ffffff",
   75418 => x"ffffff",
   75419 => x"ffffff",
   75420 => x"ffffff",
   75421 => x"ffffff",
   75422 => x"ffffff",
   75423 => x"ffffff",
   75424 => x"ffffff",
   75425 => x"ffffff",
   75426 => x"ffffff",
   75427 => x"ffffff",
   75428 => x"ffffff",
   75429 => x"ffffff",
   75430 => x"ffffff",
   75431 => x"ffffff",
   75432 => x"ffffff",
   75433 => x"ffffff",
   75434 => x"ffffff",
   75435 => x"ffffff",
   75436 => x"ffffff",
   75437 => x"ffffff",
   75438 => x"ffffff",
   75439 => x"ffffff",
   75440 => x"ffffff",
   75441 => x"ffffff",
   75442 => x"ffffff",
   75443 => x"ffffff",
   75444 => x"ffffff",
   75445 => x"ffffff",
   75446 => x"ffffff",
   75447 => x"ffffff",
   75448 => x"ffffff",
   75449 => x"ffffff",
   75450 => x"ffffff",
   75451 => x"ffffff",
   75452 => x"ffffff",
   75453 => x"ffffff",
   75454 => x"ffffff",
   75455 => x"ffffff",
   75456 => x"ffffff",
   75457 => x"ffffff",
   75458 => x"ffffff",
   75459 => x"ffffff",
   75460 => x"ffffff",
   75461 => x"ffffff",
   75462 => x"ffffff",
   75463 => x"ffffff",
   75464 => x"ffffff",
   75465 => x"ffffff",
   75466 => x"ffffff",
   75467 => x"ffffff",
   75468 => x"ffffff",
   75469 => x"ffffff",
   75470 => x"ffffff",
   75471 => x"ffffff",
   75472 => x"ffffff",
   75473 => x"ffffff",
   75474 => x"ffffff",
   75475 => x"ffffff",
   75476 => x"ffffff",
   75477 => x"ffffff",
   75478 => x"ffffff",
   75479 => x"ffffff",
   75480 => x"ffffff",
   75481 => x"ffffff",
   75482 => x"ffffff",
   75483 => x"ffffff",
   75484 => x"ffffff",
   75485 => x"ffffff",
   75486 => x"ffffff",
   75487 => x"ffffff",
   75488 => x"ffffff",
   75489 => x"ffffff",
   75490 => x"ffffff",
   75491 => x"ffffff",
   75492 => x"ffffff",
   75493 => x"ffffff",
   75494 => x"ffffff",
   75495 => x"ffffff",
   75496 => x"ffffff",
   75497 => x"ffffff",
   75498 => x"ffffff",
   75499 => x"ffffff",
   75500 => x"ffffff",
   75501 => x"ffffff",
   75502 => x"ffffff",
   75503 => x"ffffff",
   75504 => x"ffffff",
   75505 => x"ffffff",
   75506 => x"ffffff",
   75507 => x"ffffff",
   75508 => x"ffffff",
   75509 => x"ffffff",
   75510 => x"ffffff",
   75511 => x"ffffff",
   75512 => x"ffffff",
   75513 => x"ffffff",
   75514 => x"ffffff",
   75515 => x"ffffff",
   75516 => x"ffffff",
   75517 => x"ffffff",
   75518 => x"ffffff",
   75519 => x"ffffff",
   75520 => x"ffffff",
   75521 => x"ffffff",
   75522 => x"ffffff",
   75523 => x"ffffff",
   75524 => x"ffffff",
   75525 => x"ffffff",
   75526 => x"ffffff",
   75527 => x"ffffff",
   75528 => x"ffffff",
   75529 => x"ffffff",
   75530 => x"ffffff",
   75531 => x"ffffff",
   75532 => x"ffffff",
   75533 => x"ffffff",
   75534 => x"ffffff",
   75535 => x"ffffff",
   75536 => x"ffffff",
   75537 => x"ffffff",
   75538 => x"ffffff",
   75539 => x"ffffff",
   75540 => x"ffffff",
   75541 => x"ffffff",
   75542 => x"ffffff",
   75543 => x"ffffff",
   75544 => x"ffffff",
   75545 => x"ffffff",
   75546 => x"ffffff",
   75547 => x"ffffff",
   75548 => x"ffffff",
   75549 => x"ffffff",
   75550 => x"ffffff",
   75551 => x"ffffff",
   75552 => x"ffffff",
   75553 => x"ffffff",
   75554 => x"ffffff",
   75555 => x"ffffff",
   75556 => x"ffffff",
   75557 => x"ffffff",
   75558 => x"ffffff",
   75559 => x"ffffff",
   75560 => x"ffffff",
   75561 => x"ffffff",
   75562 => x"ffffff",
   75563 => x"ffffff",
   75564 => x"ffffff",
   75565 => x"ffffff",
   75566 => x"ffffff",
   75567 => x"ffffff",
   75568 => x"ffffff",
   75569 => x"ffffff",
   75570 => x"ffffff",
   75571 => x"ffffff",
   75572 => x"ffffff",
   75573 => x"ffffff",
   75574 => x"ffffff",
   75575 => x"ffffff",
   75576 => x"ffffff",
   75577 => x"ffffff",
   75578 => x"ffffff",
   75579 => x"ffffff",
   75580 => x"ffffff",
   75581 => x"ffffff",
   75582 => x"ffffff",
   75583 => x"ffffff",
   75584 => x"ffffff",
   75585 => x"ffffff",
   75586 => x"ffffff",
   75587 => x"ffffff",
   75588 => x"ffffff",
   75589 => x"ffffff",
   75590 => x"ffffff",
   75591 => x"ffffff",
   75592 => x"ffffff",
   75593 => x"ffffff",
   75594 => x"ffffff",
   75595 => x"ffffff",
   75596 => x"ffffff",
   75597 => x"ffffff",
   75598 => x"ffffff",
   75599 => x"ffffff",
   75600 => x"ffffff",
   75601 => x"ffffff",
   75602 => x"ffffff",
   75603 => x"ffffff",
   75604 => x"ffffff",
   75605 => x"ffffff",
   75606 => x"ffffff",
   75607 => x"ffffff",
   75608 => x"ffffff",
   75609 => x"ffffff",
   75610 => x"ffffff",
   75611 => x"ffffff",
   75612 => x"ffffff",
   75613 => x"ffffff",
   75614 => x"ffffff",
   75615 => x"ffffff",
   75616 => x"ffffff",
   75617 => x"ffffff",
   75618 => x"ffffff",
   75619 => x"ffffff",
   75620 => x"ffffff",
   75621 => x"ffffff",
   75622 => x"ffffff",
   75623 => x"ffffff",
   75624 => x"ffffff",
   75625 => x"ffffff",
   75626 => x"ffffff",
   75627 => x"ffffff",
   75628 => x"ffffff",
   75629 => x"ffffff",
   75630 => x"ffffff",
   75631 => x"ffffff",
   75632 => x"ffffff",
   75633 => x"ffffff",
   75634 => x"ffffff",
   75635 => x"ffffff",
   75636 => x"ffffff",
   75637 => x"ffffff",
   75638 => x"ffffff",
   75639 => x"ffffff",
   75640 => x"ffffff",
   75641 => x"ffffff",
   75642 => x"ffffff",
   75643 => x"ffffff",
   75644 => x"ffffff",
   75645 => x"ffffff",
   75646 => x"ffffff",
   75647 => x"ffffff",
   75648 => x"ffffff",
   75649 => x"ffffff",
   75650 => x"ffffff",
   75651 => x"ffffff",
   75652 => x"ffffff",
   75653 => x"ffffff",
   75654 => x"ffffff",
   75655 => x"ffffff",
   75656 => x"ffffff",
   75657 => x"ffffff",
   75658 => x"ffffff",
   75659 => x"ffffff",
   75660 => x"ffffff",
   75661 => x"ffffff",
   75662 => x"ffffff",
   75663 => x"ffffff",
   75664 => x"ffffff",
   75665 => x"ffffff",
   75666 => x"ffffff",
   75667 => x"ffffff",
   75668 => x"ffffff",
   75669 => x"ffffff",
   75670 => x"ffffff",
   75671 => x"ffffff",
   75672 => x"ffffff",
   75673 => x"ffffff",
   75674 => x"ffffff",
   75675 => x"ffffff",
   75676 => x"ffffff",
   75677 => x"ffffff",
   75678 => x"ffffff",
   75679 => x"ffffff",
   75680 => x"ffffff",
   75681 => x"ffffff",
   75682 => x"ffffff",
   75683 => x"ffffff",
   75684 => x"ffffff",
   75685 => x"ffffff",
   75686 => x"ffffff",
   75687 => x"ffffff",
   75688 => x"ffffff",
   75689 => x"ffffff",
   75690 => x"ffffff",
   75691 => x"ffffff",
   75692 => x"ffffff",
   75693 => x"ffffff",
   75694 => x"ffffff",
   75695 => x"ffffff",
   75696 => x"ffffff",
   75697 => x"ffffff",
   75698 => x"ffffff",
   75699 => x"ffffff",
   75700 => x"ffffff",
   75701 => x"ffffff",
   75702 => x"ffffff",
   75703 => x"ffffff",
   75704 => x"ffffff",
   75705 => x"ffffff",
   75706 => x"ffffff",
   75707 => x"ffffff",
   75708 => x"ffffff",
   75709 => x"ffffff",
   75710 => x"ffffff",
   75711 => x"ffffff",
   75712 => x"ffffff",
   75713 => x"ffffff",
   75714 => x"ffffff",
   75715 => x"ffffff",
   75716 => x"ffffff",
   75717 => x"ffffff",
   75718 => x"ffffff",
   75719 => x"ffffff",
   75720 => x"ffffff",
   75721 => x"ffffff",
   75722 => x"ffffff",
   75723 => x"ffffff",
   75724 => x"ffffff",
   75725 => x"ffffff",
   75726 => x"ffffff",
   75727 => x"ffffff",
   75728 => x"ffffff",
   75729 => x"ffffff",
   75730 => x"ffffff",
   75731 => x"ffffff",
   75732 => x"ffffff",
   75733 => x"ffffff",
   75734 => x"ffffff",
   75735 => x"ffffff",
   75736 => x"ffffff",
   75737 => x"ffffff",
   75738 => x"ffffff",
   75739 => x"ffffff",
   75740 => x"ffffff",
   75741 => x"ffffff",
   75742 => x"ffffff",
   75743 => x"ffffff",
   75744 => x"ffffff",
   75745 => x"ffffff",
   75746 => x"ffffff",
   75747 => x"ffffff",
   75748 => x"ffffff",
   75749 => x"ffffff",
   75750 => x"ffffff",
   75751 => x"ffffff",
   75752 => x"ffffff",
   75753 => x"ffffff",
   75754 => x"ffffff",
   75755 => x"ffffff",
   75756 => x"ffffff",
   75757 => x"ffffff",
   75758 => x"ffffff",
   75759 => x"ffffff",
   75760 => x"ffffff",
   75761 => x"ffffff",
   75762 => x"ffffff",
   75763 => x"ffffff",
   75764 => x"ffffff",
   75765 => x"ffffff",
   75766 => x"ffffff",
   75767 => x"ffffff",
   75768 => x"ffffff",
   75769 => x"ffffff",
   75770 => x"ffffff",
   75771 => x"ffffff",
   75772 => x"ffffff",
   75773 => x"ffffff",
   75774 => x"ffffff",
   75775 => x"ffffff",
   75776 => x"ffffff",
   75777 => x"ffffff",
   75778 => x"ffffff",
   75779 => x"ffffff",
   75780 => x"ffffff",
   75781 => x"ffffff",
   75782 => x"ffffff",
   75783 => x"ffffff",
   75784 => x"ffffff",
   75785 => x"ffffff",
   75786 => x"ffffff",
   75787 => x"ffffff",
   75788 => x"ffffff",
   75789 => x"ffffff",
   75790 => x"ffffff",
   75791 => x"ffffff",
   75792 => x"ffffff",
   75793 => x"ffffff",
   75794 => x"ffffff",
   75795 => x"ffffff",
   75796 => x"ffffff",
   75797 => x"ffffff",
   75798 => x"ffffff",
   75799 => x"ffffff",
   75800 => x"ffffff",
   75801 => x"ffffff",
   75802 => x"ffffff",
   75803 => x"ffffff",
   75804 => x"ffffff",
   75805 => x"ffffff",
   75806 => x"ffffff",
   75807 => x"ffffff",
   75808 => x"ffffff",
   75809 => x"ffffff",
   75810 => x"ffffff",
   75811 => x"ffffff",
   75812 => x"ffffff",
   75813 => x"ffffff",
   75814 => x"ffffff",
   75815 => x"ffffff",
   75816 => x"ffffff",
   75817 => x"ffffff",
   75818 => x"ffffff",
   75819 => x"ffffff",
   75820 => x"ffffff",
   75821 => x"ffffff",
   75822 => x"ffffff",
   75823 => x"ffffff",
   75824 => x"ffffff",
   75825 => x"ffffff",
   75826 => x"ffffff",
   75827 => x"ffffff",
   75828 => x"ffffff",
   75829 => x"ffffff",
   75830 => x"ffffff",
   75831 => x"ffffff",
   75832 => x"ffffff",
   75833 => x"ffffff",
   75834 => x"ffffff",
   75835 => x"ffffff",
   75836 => x"ffffff",
   75837 => x"ffffff",
   75838 => x"ffffff",
   75839 => x"ffffff",
   75840 => x"ffffff",
   75841 => x"ffffff",
   75842 => x"ffffff",
   75843 => x"ffffff",
   75844 => x"ffffff",
   75845 => x"ffffff",
   75846 => x"ffffff",
   75847 => x"ffffff",
   75848 => x"ffffff",
   75849 => x"ffffff",
   75850 => x"ffffff",
   75851 => x"ffffff",
   75852 => x"ffffff",
   75853 => x"ffffff",
   75854 => x"ffffff",
   75855 => x"ffffff",
   75856 => x"ffffff",
   75857 => x"ffffff",
   75858 => x"ffffff",
   75859 => x"ffffff",
   75860 => x"ffffff",
   75861 => x"ffffff",
   75862 => x"ffffff",
   75863 => x"ffffff",
   75864 => x"ffffff",
   75865 => x"ffffff",
   75866 => x"ffffff",
   75867 => x"ffffff",
   75868 => x"ffffff",
   75869 => x"ffffff",
   75870 => x"ffffff",
   75871 => x"ffffff",
   75872 => x"ffffff",
   75873 => x"ffffff",
   75874 => x"ffffff",
   75875 => x"ffffff",
   75876 => x"ffffff",
   75877 => x"ffffff",
   75878 => x"ffffff",
   75879 => x"ffffff",
   75880 => x"ffffff",
   75881 => x"ffffff",
   75882 => x"ffffff",
   75883 => x"ffffff",
   75884 => x"ffffff",
   75885 => x"ffffff",
   75886 => x"ffffff",
   75887 => x"ffffff",
   75888 => x"ffffff",
   75889 => x"ffffff",
   75890 => x"ffffff",
   75891 => x"ffffff",
   75892 => x"ffffff",
   75893 => x"ffffff",
   75894 => x"ffffff",
   75895 => x"ffffff",
   75896 => x"ffffff",
   75897 => x"ffffff",
   75898 => x"ffffff",
   75899 => x"ffffff",
   75900 => x"ffffff",
   75901 => x"ffffff",
   75902 => x"ffffff",
   75903 => x"ffffff",
   75904 => x"ffffff",
   75905 => x"ffffff",
   75906 => x"ffffff",
   75907 => x"ffffff",
   75908 => x"ffffff",
   75909 => x"ffffff",
   75910 => x"ffffff",
   75911 => x"ffffff",
   75912 => x"ffffff",
   75913 => x"ffffff",
   75914 => x"ffffff",
   75915 => x"ffffff",
   75916 => x"ffffff",
   75917 => x"ffffff",
   75918 => x"ffffff",
   75919 => x"ffffff",
   75920 => x"ffffff",
   75921 => x"ffffff",
   75922 => x"ffffff",
   75923 => x"ffffff",
   75924 => x"ffffff",
   75925 => x"ffffff",
   75926 => x"ffffff",
   75927 => x"ffffff",
   75928 => x"ffffff",
   75929 => x"ffffff",
   75930 => x"ffffff",
   75931 => x"ffffff",
   75932 => x"ffffff",
   75933 => x"ffffff",
   75934 => x"ffffff",
   75935 => x"ffffff",
   75936 => x"ffffff",
   75937 => x"ffffff",
   75938 => x"ffffff",
   75939 => x"ffffff",
   75940 => x"ffffff",
   75941 => x"ffffff",
   75942 => x"ffffff",
   75943 => x"ffffff",
   75944 => x"ffffff",
   75945 => x"ffffff",
   75946 => x"ffffff",
   75947 => x"ffffff",
   75948 => x"ffffff",
   75949 => x"ffffff",
   75950 => x"ffffff",
   75951 => x"ffffff",
   75952 => x"ffffff",
   75953 => x"ffffff",
   75954 => x"ffffff",
   75955 => x"ffffff",
   75956 => x"ffffff",
   75957 => x"ffffff",
   75958 => x"ffffff",
   75959 => x"ffffff",
   75960 => x"ffffff",
   75961 => x"ffffff",
   75962 => x"ffffff",
   75963 => x"ffffff",
   75964 => x"ffffff",
   75965 => x"ffffff",
   75966 => x"ffffff",
   75967 => x"ffffff",
   75968 => x"ffffff",
   75969 => x"ffffff",
   75970 => x"ffffff",
   75971 => x"ffffff",
   75972 => x"ffffff",
   75973 => x"ffffff",
   75974 => x"ffffff",
   75975 => x"ffffff",
   75976 => x"ffffff",
   75977 => x"ffffff",
   75978 => x"ffffff",
   75979 => x"ffffff",
   75980 => x"ffffff",
   75981 => x"ffffff",
   75982 => x"ffffff",
   75983 => x"ffffff",
   75984 => x"ffffff",
   75985 => x"ffffff",
   75986 => x"ffffff",
   75987 => x"ffffff",
   75988 => x"ffffff",
   75989 => x"ffffff",
   75990 => x"ffffff",
   75991 => x"ffffff",
   75992 => x"ffffff",
   75993 => x"ffffff",
   75994 => x"ffffff",
   75995 => x"ffffff",
   75996 => x"ffffff",
   75997 => x"ffffff",
   75998 => x"ffffff",
   75999 => x"ffffff",
   76000 => x"ffffff",
   76001 => x"ffffff",
   76002 => x"ffffff",
   76003 => x"ffffff",
   76004 => x"ffffff",
   76005 => x"ffffff",
   76006 => x"ffffff",
   76007 => x"ffffff",
   76008 => x"ffffff",
   76009 => x"ffffff",
   76010 => x"ffffff",
   76011 => x"ffffff",
   76012 => x"ffffff",
   76013 => x"ffffff",
   76014 => x"ffffff",
   76015 => x"ffffff",
   76016 => x"ffffff",
   76017 => x"ffffff",
   76018 => x"ffffff",
   76019 => x"ffffff",
   76020 => x"ffffff",
   76021 => x"ffffff",
   76022 => x"ffffff",
   76023 => x"ffffff",
   76024 => x"ffffff",
   76025 => x"ffffff",
   76026 => x"ffffff",
   76027 => x"ffffff",
   76028 => x"ffffff",
   76029 => x"ffffff",
   76030 => x"ffffff",
   76031 => x"ffffff",
   76032 => x"ffffff",
   76033 => x"ffffff",
   76034 => x"ffffff",
   76035 => x"ffffff",
   76036 => x"ffffff",
   76037 => x"ffffff",
   76038 => x"ffffff",
   76039 => x"ffffff",
   76040 => x"ffffff",
   76041 => x"ffffff",
   76042 => x"ffffff",
   76043 => x"ffffff",
   76044 => x"ffffff",
   76045 => x"ffffff",
   76046 => x"ffffff",
   76047 => x"ffffff",
   76048 => x"ffffff",
   76049 => x"ffffff",
   76050 => x"ffffff",
   76051 => x"ffffff",
   76052 => x"ffffff",
   76053 => x"ffffff",
   76054 => x"ffffff",
   76055 => x"ffffff",
   76056 => x"ffffff",
   76057 => x"ffffff",
   76058 => x"ffffff",
   76059 => x"ffffff",
   76060 => x"ffffff",
   76061 => x"ffffff",
   76062 => x"ffffff",
   76063 => x"ffffff",
   76064 => x"ffffff",
   76065 => x"ffffff",
   76066 => x"ffffff",
   76067 => x"ffffff",
   76068 => x"ffffff",
   76069 => x"ffffff",
   76070 => x"ffffff",
   76071 => x"ffffff",
   76072 => x"ffffff",
   76073 => x"ffffff",
   76074 => x"ffffff",
   76075 => x"ffffff",
   76076 => x"ffffff",
   76077 => x"ffffff",
   76078 => x"ffffff",
   76079 => x"ffffff",
   76080 => x"ffffff",
   76081 => x"ffffff",
   76082 => x"ffffff",
   76083 => x"ffffff",
   76084 => x"ffffff",
   76085 => x"ffffff",
   76086 => x"ffffff",
   76087 => x"ffffff",
   76088 => x"ffffff",
   76089 => x"ffffff",
   76090 => x"ffffff",
   76091 => x"ffffff",
   76092 => x"ffffff",
   76093 => x"ffffff",
   76094 => x"ffffff",
   76095 => x"ffffff",
   76096 => x"ffffff",
   76097 => x"ffffff",
   76098 => x"ffffff",
   76099 => x"ffffff",
   76100 => x"ffffff",
   76101 => x"ffffff",
   76102 => x"ffffff",
   76103 => x"ffffff",
   76104 => x"ffffff",
   76105 => x"ffffff",
   76106 => x"ffffff",
   76107 => x"ffffff",
   76108 => x"ffffff",
   76109 => x"ffffff",
   76110 => x"ffffff",
   76111 => x"ffffff",
   76112 => x"ffffff",
   76113 => x"ffffff",
   76114 => x"ffffff",
   76115 => x"ffffff",
   76116 => x"ffffff",
   76117 => x"ffffff",
   76118 => x"ffffff",
   76119 => x"ffffff",
   76120 => x"ffffff",
   76121 => x"ffffff",
   76122 => x"ffffff",
   76123 => x"ffffff",
   76124 => x"ffffff",
   76125 => x"ffffff",
   76126 => x"ffffff",
   76127 => x"ffffff",
   76128 => x"ffffff",
   76129 => x"ffffff",
   76130 => x"ffffff",
   76131 => x"ffffff",
   76132 => x"ffffff",
   76133 => x"ffffff",
   76134 => x"ffffff",
   76135 => x"ffffff",
   76136 => x"ffffff",
   76137 => x"ffffff",
   76138 => x"ffffff",
   76139 => x"ffffff",
   76140 => x"ffffff",
   76141 => x"ffffff",
   76142 => x"ffffff",
   76143 => x"ffffff",
   76144 => x"ffffff",
   76145 => x"ffffff",
   76146 => x"ffffff",
   76147 => x"ffffff",
   76148 => x"ffffff",
   76149 => x"ffffff",
   76150 => x"ffffff",
   76151 => x"ffffff",
   76152 => x"ffffff",
   76153 => x"ffffff",
   76154 => x"ffffff",
   76155 => x"ffffff",
   76156 => x"ffffff",
   76157 => x"ffffff",
   76158 => x"ffffff",
   76159 => x"ffffff",
   76160 => x"ffffff",
   76161 => x"ffffff",
   76162 => x"ffffff",
   76163 => x"ffffff",
   76164 => x"ffffff",
   76165 => x"ffffff",
   76166 => x"ffffff",
   76167 => x"ffffff",
   76168 => x"ffffff",
   76169 => x"ffffff",
   76170 => x"ffffff",
   76171 => x"ffffff",
   76172 => x"ffffff",
   76173 => x"ffffff",
   76174 => x"ffffff",
   76175 => x"ffffff",
   76176 => x"ffffff",
   76177 => x"ffffff",
   76178 => x"ffffff",
   76179 => x"ffffff",
   76180 => x"ffffff",
   76181 => x"ffffff",
   76182 => x"ffffff",
   76183 => x"ffffff",
   76184 => x"ffffff",
   76185 => x"ffffff",
   76186 => x"ffffff",
   76187 => x"ffffff",
   76188 => x"ffffff",
   76189 => x"ffffff",
   76190 => x"ffffff",
   76191 => x"ffffff",
   76192 => x"ffffff",
   76193 => x"ffffff",
   76194 => x"ffffff",
   76195 => x"ffffff",
   76196 => x"ffffff",
   76197 => x"ffffff",
   76198 => x"ffffff",
   76199 => x"ffffff",
   76200 => x"ffffff",
   76201 => x"ffffff",
   76202 => x"ffffff",
   76203 => x"ffffff",
   76204 => x"ffffff",
   76205 => x"ffffff",
   76206 => x"ffffff",
   76207 => x"ffffff",
   76208 => x"ffffff",
   76209 => x"ffffff",
   76210 => x"ffffff",
   76211 => x"ffffff",
   76212 => x"ffffff",
   76213 => x"ffffff",
   76214 => x"ffffff",
   76215 => x"ffffff",
   76216 => x"ffffff",
   76217 => x"ffffff",
   76218 => x"ffffff",
   76219 => x"ffffff",
   76220 => x"ffffff",
   76221 => x"ffffff",
   76222 => x"ffffff",
   76223 => x"ffffff",
   76224 => x"ffffff",
   76225 => x"ffffff",
   76226 => x"ffffff",
   76227 => x"ffffff",
   76228 => x"ffffff",
   76229 => x"ffffff",
   76230 => x"ffffff",
   76231 => x"ffffff",
   76232 => x"ffffff",
   76233 => x"ffffff",
   76234 => x"ffffff",
   76235 => x"ffffff",
   76236 => x"ffffff",
   76237 => x"ffffff",
   76238 => x"ffffff",
   76239 => x"ffffff",
   76240 => x"ffffff",
   76241 => x"ffffff",
   76242 => x"ffffff",
   76243 => x"ffffff",
   76244 => x"ffffff",
   76245 => x"ffffff",
   76246 => x"ffffff",
   76247 => x"ffffff",
   76248 => x"ffffff",
   76249 => x"ffffff",
   76250 => x"ffffff",
   76251 => x"ffffff",
   76252 => x"ffffff",
   76253 => x"ffffff",
   76254 => x"ffffff",
   76255 => x"ffffff",
   76256 => x"ffffff",
   76257 => x"ffffff",
   76258 => x"ffffff",
   76259 => x"ffffff",
   76260 => x"ffffff",
   76261 => x"ffffff",
   76262 => x"ffffff",
   76263 => x"ffffff",
   76264 => x"ffffff",
   76265 => x"ffffff",
   76266 => x"ffffff",
   76267 => x"ffffff",
   76268 => x"ffffff",
   76269 => x"ffffff",
   76270 => x"ffffff",
   76271 => x"ffffff",
   76272 => x"ffffff",
   76273 => x"ffffff",
   76274 => x"ffffff",
   76275 => x"ffffff",
   76276 => x"ffffff",
   76277 => x"ffffff",
   76278 => x"ffffff",
   76279 => x"ffffff",
   76280 => x"ffffff",
   76281 => x"ffffff",
   76282 => x"ffffff",
   76283 => x"ffffff",
   76284 => x"ffffff",
   76285 => x"ffffff",
   76286 => x"ffffff",
   76287 => x"ffffff",
   76288 => x"ffffff",
   76289 => x"ffffff",
   76290 => x"ffffff",
   76291 => x"ffffff",
   76292 => x"ffffff",
   76293 => x"ffffff",
   76294 => x"ffffff",
   76295 => x"ffffff",
   76296 => x"ffffff",
   76297 => x"ffffff",
   76298 => x"ffffff",
   76299 => x"ffffff",
   76300 => x"ffffff",
   76301 => x"ffffff",
   76302 => x"ffffff",
   76303 => x"ffffff",
   76304 => x"ffffff",
   76305 => x"ffffff",
   76306 => x"ffffff",
   76307 => x"ffffff",
   76308 => x"ffffff",
   76309 => x"ffffff",
   76310 => x"ffffff",
   76311 => x"ffffff",
   76312 => x"ffffff",
   76313 => x"ffffff",
   76314 => x"ffffff",
   76315 => x"ffffff",
   76316 => x"ffffff",
   76317 => x"ffffff",
   76318 => x"ffffff",
   76319 => x"ffffff",
   76320 => x"ffffff",
   76321 => x"ffffff",
   76322 => x"ffffff",
   76323 => x"ffffff",
   76324 => x"ffffff",
   76325 => x"ffffff",
   76326 => x"ffffff",
   76327 => x"ffffff",
   76328 => x"ffffff",
   76329 => x"ffffff",
   76330 => x"ffffff",
   76331 => x"ffffff",
   76332 => x"ffffff",
   76333 => x"ffffff",
   76334 => x"ffffff",
   76335 => x"ffffff",
   76336 => x"ffffff",
   76337 => x"ffffff",
   76338 => x"ffffff",
   76339 => x"ffffff",
   76340 => x"ffffff",
   76341 => x"ffffff",
   76342 => x"ffffff",
   76343 => x"ffffff",
   76344 => x"ffffff",
   76345 => x"ffffff",
   76346 => x"ffffff",
   76347 => x"ffffff",
   76348 => x"ffffff",
   76349 => x"ffffff",
   76350 => x"ffffff",
   76351 => x"ffffff",
   76352 => x"ffffff",
   76353 => x"ffffff",
   76354 => x"ffffff",
   76355 => x"ffffff",
   76356 => x"ffffff",
   76357 => x"ffffff",
   76358 => x"ffffff",
   76359 => x"ffffff",
   76360 => x"ffffff",
   76361 => x"ffffff",
   76362 => x"ffffff",
   76363 => x"ffffff",
   76364 => x"ffffff",
   76365 => x"ffffff",
   76366 => x"ffffff",
   76367 => x"ffffff",
   76368 => x"ffffff",
   76369 => x"ffffff",
   76370 => x"ffffff",
   76371 => x"ffffff",
   76372 => x"ffffff",
   76373 => x"ffffff",
   76374 => x"ffffff",
   76375 => x"ffffff",
   76376 => x"ffffff",
   76377 => x"ffffff",
   76378 => x"ffffff",
   76379 => x"ffffff",
   76380 => x"ffffff",
   76381 => x"ffffff",
   76382 => x"ffffff",
   76383 => x"ffffff",
   76384 => x"ffffff",
   76385 => x"ffffff",
   76386 => x"ffffff",
   76387 => x"ffffff",
   76388 => x"ffffff",
   76389 => x"ffffff",
   76390 => x"ffffff",
   76391 => x"ffffff",
   76392 => x"ffffff",
   76393 => x"ffffff",
   76394 => x"ffffff",
   76395 => x"ffffff",
   76396 => x"ffffff",
   76397 => x"ffffff",
   76398 => x"ffffff",
   76399 => x"ffffff",
   76400 => x"ffffff",
   76401 => x"ffffff",
   76402 => x"ffffff",
   76403 => x"ffffff",
   76404 => x"ffffff",
   76405 => x"ffffff",
   76406 => x"ffffff",
   76407 => x"ffffff",
   76408 => x"ffffff",
   76409 => x"ffffff",
   76410 => x"ffffff",
   76411 => x"ffffff",
   76412 => x"ffffff",
   76413 => x"ffffff",
   76414 => x"ffffff",
   76415 => x"ffffff",
   76416 => x"ffffff",
   76417 => x"ffffff",
   76418 => x"ffffff",
   76419 => x"ffffff",
   76420 => x"ffffff",
   76421 => x"ffffff",
   76422 => x"ffffff",
   76423 => x"ffffff",
   76424 => x"ffffff",
   76425 => x"ffffff",
   76426 => x"ffffff",
   76427 => x"ffffff",
   76428 => x"ffffff",
   76429 => x"ffffff",
   76430 => x"ffffff",
   76431 => x"ffffff",
   76432 => x"ffffff",
   76433 => x"ffffff",
   76434 => x"ffffff",
   76435 => x"ffffff",
   76436 => x"ffffff",
   76437 => x"ffffff",
   76438 => x"ffffff",
   76439 => x"ffffff",
   76440 => x"ffffff",
   76441 => x"ffffff",
   76442 => x"ffffff",
   76443 => x"ffffff",
   76444 => x"ffffff",
   76445 => x"ffffff",
   76446 => x"ffffff",
   76447 => x"ffffff",
   76448 => x"ffffff",
   76449 => x"ffffff",
   76450 => x"ffffff",
   76451 => x"ffffff",
   76452 => x"ffffff",
   76453 => x"ffffff",
   76454 => x"ffffff",
   76455 => x"ffffff",
   76456 => x"ffffff",
   76457 => x"ffffff",
   76458 => x"ffffff",
   76459 => x"ffffff",
   76460 => x"ffffff",
   76461 => x"ffffff",
   76462 => x"ffffff",
   76463 => x"ffffff",
   76464 => x"ffffff",
   76465 => x"ffffff",
   76466 => x"ffffff",
   76467 => x"ffffff",
   76468 => x"ffffff",
   76469 => x"ffffff",
   76470 => x"ffffff",
   76471 => x"ffffff",
   76472 => x"ffffff",
   76473 => x"ffffff",
   76474 => x"ffffff",
   76475 => x"ffffff",
   76476 => x"ffffff",
   76477 => x"ffffff",
   76478 => x"ffffff",
   76479 => x"ffffff",
   76480 => x"ffffff",
   76481 => x"ffffff",
   76482 => x"ffffff",
   76483 => x"ffffff",
   76484 => x"ffffff",
   76485 => x"ffffff",
   76486 => x"ffffff",
   76487 => x"ffffff",
   76488 => x"ffffff",
   76489 => x"ffffff",
   76490 => x"ffffff",
   76491 => x"ffffff",
   76492 => x"ffffff",
   76493 => x"ffffff",
   76494 => x"ffffff",
   76495 => x"ffffff",
   76496 => x"ffffff",
   76497 => x"ffffff",
   76498 => x"ffffff",
   76499 => x"ffffff",
   76500 => x"ffffff",
   76501 => x"ffffff",
   76502 => x"ffffff",
   76503 => x"ffffff",
   76504 => x"ffffff",
   76505 => x"ffffff",
   76506 => x"ffffff",
   76507 => x"ffffff",
   76508 => x"ffffff",
   76509 => x"ffffff",
   76510 => x"ffffff",
   76511 => x"ffffff",
   76512 => x"ffffff",
   76513 => x"ffffff",
   76514 => x"ffffff",
   76515 => x"ffffff",
   76516 => x"ffffff",
   76517 => x"ffffff",
   76518 => x"ffffff",
   76519 => x"ffffff",
   76520 => x"ffffff",
   76521 => x"ffffff",
   76522 => x"ffffff",
   76523 => x"ffffff",
   76524 => x"ffffff",
   76525 => x"ffffff",
   76526 => x"ffffff",
   76527 => x"ffffff",
   76528 => x"ffffff",
   76529 => x"ffffff",
   76530 => x"ffffff",
   76531 => x"ffffff",
   76532 => x"ffffff",
   76533 => x"ffffff",
   76534 => x"ffffff",
   76535 => x"ffffff",
   76536 => x"ffffff",
   76537 => x"ffffff",
   76538 => x"ffffff",
   76539 => x"ffffff",
   76540 => x"ffffff",
   76541 => x"ffffff",
   76542 => x"ffffff",
   76543 => x"ffffff",
   76544 => x"ffffff",
   76545 => x"ffffff",
   76546 => x"ffffff",
   76547 => x"ffffff",
   76548 => x"ffffff",
   76549 => x"ffffff",
   76550 => x"ffffff",
   76551 => x"ffffff",
   76552 => x"ffffff",
   76553 => x"ffffff",
   76554 => x"ffffff",
   76555 => x"ffffff",
   76556 => x"ffffff",
   76557 => x"ffffff",
   76558 => x"ffffff",
   76559 => x"ffffff",
   76560 => x"ffffff",
   76561 => x"ffffff",
   76562 => x"ffffff",
   76563 => x"ffffff",
   76564 => x"ffffff",
   76565 => x"ffffff",
   76566 => x"ffffff",
   76567 => x"ffffff",
   76568 => x"ffffff",
   76569 => x"ffffff",
   76570 => x"ffffff",
   76571 => x"ffffff",
   76572 => x"ffffff",
   76573 => x"ffffff",
   76574 => x"ffffff",
   76575 => x"ffffff",
   76576 => x"ffffff",
   76577 => x"ffffff",
   76578 => x"ffffff",
   76579 => x"ffffff",
   76580 => x"ffffff",
   76581 => x"ffffff",
   76582 => x"ffffff",
   76583 => x"ffffff",
   76584 => x"ffffff",
   76585 => x"ffffff",
   76586 => x"ffffff",
   76587 => x"ffffff",
   76588 => x"ffffff",
   76589 => x"ffffff",
   76590 => x"ffffff",
   76591 => x"ffffff",
   76592 => x"ffffff",
   76593 => x"ffffff",
   76594 => x"ffffff",
   76595 => x"ffffff",
   76596 => x"ffffff",
   76597 => x"ffffff",
   76598 => x"ffffff",
   76599 => x"ffffff",
   76600 => x"ffffff",
   76601 => x"ffffff",
   76602 => x"ffffff",
   76603 => x"ffffff",
   76604 => x"ffffff",
   76605 => x"ffffff",
   76606 => x"ffffff",
   76607 => x"ffffff",
   76608 => x"ffffff",
   76609 => x"ffffff",
   76610 => x"ffffff",
   76611 => x"ffffff",
   76612 => x"ffffff",
   76613 => x"ffffff",
   76614 => x"ffffff",
   76615 => x"ffffff",
   76616 => x"ffffff",
   76617 => x"ffffff",
   76618 => x"ffffff",
   76619 => x"ffffff",
   76620 => x"ffffff",
   76621 => x"ffffff",
   76622 => x"ffffff",
   76623 => x"ffffff",
   76624 => x"ffffff",
   76625 => x"ffffff",
   76626 => x"ffffff",
   76627 => x"ffffff",
   76628 => x"ffffff",
   76629 => x"ffffff",
   76630 => x"ffffff",
   76631 => x"ffffff",
   76632 => x"ffffff",
   76633 => x"ffffff",
   76634 => x"ffffff",
   76635 => x"ffffff",
   76636 => x"ffffff",
   76637 => x"ffffff",
   76638 => x"ffffff",
   76639 => x"ffffff",
   76640 => x"ffffff",
   76641 => x"ffffff",
   76642 => x"ffffff",
   76643 => x"ffffff",
   76644 => x"ffffff",
   76645 => x"ffffff",
   76646 => x"ffffff",
   76647 => x"ffffff",
   76648 => x"ffffff",
   76649 => x"ffffff",
   76650 => x"ffffff",
   76651 => x"ffffff",
   76652 => x"ffffff",
   76653 => x"ffffff",
   76654 => x"ffffff",
   76655 => x"ffffff",
   76656 => x"ffffff",
   76657 => x"ffffff",
   76658 => x"ffffff",
   76659 => x"ffffff",
   76660 => x"ffffff",
   76661 => x"ffffff",
   76662 => x"ffffff",
   76663 => x"ffffff",
   76664 => x"ffffff",
   76665 => x"ffffff",
   76666 => x"ffffff",
   76667 => x"ffffff",
   76668 => x"ffffff",
   76669 => x"ffffff",
   76670 => x"ffffff",
   76671 => x"ffffff",
   76672 => x"ffffff",
   76673 => x"ffffff",
   76674 => x"ffffff",
   76675 => x"ffffff",
   76676 => x"ffffff",
   76677 => x"ffffff",
   76678 => x"ffffff",
   76679 => x"ffffff",
   76680 => x"ffffff",
   76681 => x"ffffff",
   76682 => x"ffffff",
   76683 => x"ffffff",
   76684 => x"ffffff",
   76685 => x"ffffff",
   76686 => x"ffffff",
   76687 => x"ffffff",
   76688 => x"ffffff",
   76689 => x"ffffff",
   76690 => x"ffffff",
   76691 => x"ffffff",
   76692 => x"ffffff",
   76693 => x"ffffff",
   76694 => x"ffffff",
   76695 => x"ffffff",
   76696 => x"ffffff",
   76697 => x"ffffff",
   76698 => x"ffffff",
   76699 => x"ffffff",
   76700 => x"ffffff",
   76701 => x"ffffff",
   76702 => x"ffffff",
   76703 => x"ffffff",
   76704 => x"ffffff",
   76705 => x"ffffff",
   76706 => x"ffffff",
   76707 => x"ffffff",
   76708 => x"ffffff",
   76709 => x"ffffff",
   76710 => x"ffffff",
   76711 => x"ffffff",
   76712 => x"ffffff",
   76713 => x"ffffff",
   76714 => x"ffffff",
   76715 => x"ffffff",
   76716 => x"ffffff",
   76717 => x"ffffff",
   76718 => x"ffffff",
   76719 => x"ffffff",
   76720 => x"ffffff",
   76721 => x"ffffff",
   76722 => x"ffffff",
   76723 => x"ffffff",
   76724 => x"ffffff",
   76725 => x"ffffff",
   76726 => x"ffffff",
   76727 => x"ffffff",
   76728 => x"ffffff",
   76729 => x"ffffff",
   76730 => x"ffffff",
   76731 => x"ffffff",
   76732 => x"ffffff",
   76733 => x"ffffff",
   76734 => x"ffffff",
   76735 => x"ffffff",
   76736 => x"ffffff",
   76737 => x"ffffff",
   76738 => x"ffffff",
   76739 => x"ffffff",
   76740 => x"ffffff",
   76741 => x"ffffff",
   76742 => x"ffffff",
   76743 => x"ffffff",
   76744 => x"ffffff",
   76745 => x"ffffff",
   76746 => x"ffffff",
   76747 => x"ffffff",
   76748 => x"ffffff",
   76749 => x"ffffff",
   76750 => x"ffffff",
   76751 => x"ffffff",
   76752 => x"ffffff",
   76753 => x"ffffff",
   76754 => x"ffffff",
   76755 => x"ffffff",
   76756 => x"ffffff",
   76757 => x"ffffff",
   76758 => x"ffffff",
   76759 => x"ffffff",
   76760 => x"ffffff",
   76761 => x"ffffff",
   76762 => x"ffffff",
   76763 => x"ffffff",
   76764 => x"ffffff",
   76765 => x"ffffff",
   76766 => x"ffffff",
   76767 => x"ffffff",
   76768 => x"ffffff",
   76769 => x"ffffff",
   76770 => x"ffffff",
   76771 => x"ffffff",
   76772 => x"ffffff",
   76773 => x"ffffff",
   76774 => x"ffffff",
   76775 => x"ffffff",
   76776 => x"ffffff",
   76777 => x"ffffff",
   76778 => x"ffffff",
   76779 => x"ffffff",
   76780 => x"ffffff",
   76781 => x"ffffff",
   76782 => x"ffffff",
   76783 => x"ffffff",
   76784 => x"ffffff",
   76785 => x"ffffff",
   76786 => x"ffffff",
   76787 => x"ffffff",
   76788 => x"ffffff",
   76789 => x"ffffff",
   76790 => x"ffffff",
   76791 => x"ffffff",
   76792 => x"ffffff",
   76793 => x"ffffff",
   76794 => x"ffffff",
   76795 => x"ffffff",
   76796 => x"ffffff",
   76797 => x"ffffff",
   76798 => x"ffffff",
   76799 => x"ffffff",
 others => x"FFFFFF"
    );
begin
  process(CLK)
  begin 
    if (CLK'event AND CLK='1') then
      do <= ROM(to_integer(addr));
    end if;
  end process;
end Behavioral;
