library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
use UNISIM.Vcomponents.ALL;
use work.prog_data_pkg.all;

entity RAM_VIDEO is
  port ( 
    clk  : in    std_logic;   
    addr : in    unsigned (16 downto 0); 
    do   : out   unsigned(23 downto 0);
    we   : in    std_logic
    );
end RAM_VIDEO;

architecture Behavioral of RAM_VIDEO is
  
   signal en : unsigned(37 downto 0);
   subtype mot is std_logic_vector(23 downto 0);
   type vec is array (natural range 0 to 37) of mot;
   signal DOvec : vec;
begin
        process (addr(16 downto 11),DOvec)
                variable i : integer;
        begin
                en <= (others => '0');
                i:=to_integer(addr(16 downto 11));
                en(i) <= '1';
                DO <= unsigned(DOvec(i));
        end process; 

RAM0_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM0_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM0_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM0_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM0_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM0_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM0_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM0_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM0_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM0_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM0_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM0_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM0_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM0_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM0_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM0_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM0_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM0_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM0_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM0_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM0_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM0_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM0_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM0_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM0_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM0_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM0_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM0_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM0_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM0_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM0_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM0_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM0_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM0_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM0_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM0_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM0_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM0_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM0_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM0_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM0_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM0_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM0_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM0_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM0_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM0_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM0_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM0_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM0_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM0_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM0_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM0_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM0_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM0_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM0_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM0_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM0_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM0_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM0_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM0_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM0_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM0_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM0_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM0_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM0_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(0), SSR=>'0', WE=>we, DO=>DOvec(0)(7 downto 0), DOP=>open);
RAM0_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM0_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM0_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM0_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM0_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM0_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM0_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM0_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM0_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM0_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM0_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM0_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM0_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM0_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM0_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM0_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM0_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM0_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM0_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM0_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM0_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM0_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM0_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM0_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM0_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM0_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM0_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM0_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM0_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM0_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM0_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM0_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM0_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM0_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM0_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM0_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM0_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM0_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM0_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM0_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM0_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM0_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM0_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM0_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM0_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM0_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM0_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM0_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM0_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM0_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM0_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM0_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM0_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM0_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM0_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM0_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM0_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM0_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM0_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM0_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM0_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM0_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM0_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM0_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM0_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(0), SSR=>'0', WE=>we, DO=>DOvec(0)(15 downto 8), DOP=>open);
RAM0_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM0_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM0_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM0_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM0_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM0_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM0_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM0_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM0_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM0_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM0_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM0_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM0_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM0_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM0_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM0_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM0_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM0_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM0_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM0_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM0_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM0_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM0_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM0_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM0_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM0_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM0_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM0_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM0_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM0_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM0_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM0_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM0_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM0_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM0_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM0_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM0_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM0_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM0_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM0_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM0_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM0_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM0_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM0_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM0_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM0_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM0_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM0_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM0_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM0_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM0_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM0_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM0_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM0_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM0_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM0_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM0_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM0_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM0_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM0_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM0_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM0_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM0_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM0_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM0_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(0), SSR=>'0', WE=>we, DO=>DOvec(0)(23 downto 16), DOP=>open);


RAM1_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM1_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM1_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM1_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM1_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM1_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM1_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM1_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM1_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM1_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM1_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM1_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM1_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM1_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM1_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM1_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM1_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM1_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM1_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM1_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM1_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM1_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM1_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM1_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM1_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM1_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM1_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM1_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM1_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM1_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM1_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM1_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM1_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM1_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM1_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM1_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM1_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM1_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM1_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM1_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM1_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM1_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM1_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM1_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM1_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM1_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM1_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM1_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM1_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM1_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM1_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM1_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM1_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM1_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM1_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM1_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM1_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM1_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM1_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM1_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM1_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM1_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM1_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM1_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM1_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(1), SSR=>'0', WE=>we, DO=>DOvec(1)(7 downto 0), DOP=>open);
RAM1_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM1_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM1_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM1_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM1_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM1_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM1_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM1_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM1_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM1_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM1_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM1_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM1_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM1_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM1_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM1_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM1_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM1_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM1_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM1_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM1_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM1_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM1_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM1_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM1_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM1_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM1_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM1_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM1_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM1_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM1_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM1_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM1_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM1_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM1_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM1_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM1_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM1_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM1_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM1_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM1_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM1_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM1_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM1_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM1_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM1_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM1_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM1_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM1_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM1_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM1_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM1_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM1_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM1_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM1_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM1_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM1_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM1_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM1_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM1_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM1_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM1_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM1_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM1_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM1_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(1), SSR=>'0', WE=>we, DO=>DOvec(1)(15 downto 8), DOP=>open);
RAM1_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM1_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM1_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM1_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM1_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM1_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM1_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM1_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM1_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM1_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM1_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM1_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM1_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM1_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM1_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM1_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM1_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM1_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM1_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM1_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM1_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM1_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM1_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM1_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM1_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM1_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM1_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM1_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM1_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM1_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM1_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM1_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM1_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM1_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM1_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM1_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM1_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM1_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM1_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM1_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM1_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM1_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM1_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM1_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM1_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM1_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM1_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM1_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM1_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM1_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM1_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM1_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM1_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM1_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM1_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM1_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM1_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM1_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM1_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM1_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM1_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM1_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM1_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM1_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM1_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(1), SSR=>'0', WE=>we, DO=>DOvec(1)(23 downto 16), DOP=>open);


RAM2_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM2_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM2_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM2_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM2_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM2_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM2_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM2_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM2_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM2_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM2_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM2_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM2_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM2_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM2_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM2_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM2_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM2_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM2_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM2_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM2_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM2_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM2_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM2_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM2_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM2_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM2_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM2_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM2_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM2_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM2_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM2_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM2_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM2_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM2_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM2_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM2_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM2_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM2_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM2_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM2_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM2_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM2_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM2_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM2_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM2_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM2_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM2_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM2_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM2_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM2_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM2_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM2_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM2_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM2_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM2_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM2_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM2_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM2_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM2_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM2_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM2_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM2_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM2_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM2_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(2), SSR=>'0', WE=>we, DO=>DOvec(2)(7 downto 0), DOP=>open);
RAM2_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM2_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM2_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM2_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM2_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM2_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM2_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM2_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM2_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM2_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM2_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM2_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM2_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM2_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM2_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM2_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM2_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM2_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM2_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM2_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM2_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM2_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM2_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM2_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM2_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM2_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM2_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM2_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM2_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM2_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM2_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM2_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM2_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM2_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM2_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM2_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM2_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM2_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM2_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM2_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM2_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM2_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM2_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM2_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM2_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM2_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM2_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM2_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM2_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM2_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM2_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM2_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM2_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM2_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM2_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM2_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM2_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM2_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM2_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM2_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM2_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM2_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM2_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM2_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM2_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(2), SSR=>'0', WE=>we, DO=>DOvec(2)(15 downto 8), DOP=>open);
RAM2_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM2_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM2_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM2_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM2_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM2_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM2_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM2_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM2_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM2_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM2_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM2_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM2_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM2_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM2_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM2_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM2_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM2_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM2_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM2_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM2_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM2_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM2_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM2_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM2_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM2_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM2_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM2_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM2_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM2_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM2_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM2_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM2_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM2_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM2_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM2_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM2_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM2_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM2_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM2_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM2_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM2_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM2_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM2_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM2_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM2_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM2_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM2_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM2_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM2_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM2_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM2_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM2_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM2_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM2_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM2_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM2_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM2_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM2_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM2_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM2_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM2_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM2_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM2_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM2_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(2), SSR=>'0', WE=>we, DO=>DOvec(2)(23 downto 16), DOP=>open);


RAM3_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM3_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM3_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM3_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM3_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM3_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM3_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM3_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM3_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM3_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM3_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM3_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM3_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM3_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM3_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM3_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM3_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM3_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM3_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM3_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM3_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM3_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM3_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM3_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM3_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM3_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM3_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM3_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM3_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM3_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM3_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM3_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM3_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM3_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM3_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM3_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM3_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM3_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM3_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM3_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM3_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM3_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM3_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM3_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM3_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM3_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM3_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM3_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM3_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM3_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM3_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM3_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM3_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM3_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM3_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM3_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM3_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM3_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM3_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM3_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM3_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM3_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM3_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM3_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM3_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(3), SSR=>'0', WE=>we, DO=>DOvec(3)(7 downto 0), DOP=>open);
RAM3_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM3_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM3_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM3_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM3_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM3_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM3_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM3_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM3_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM3_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM3_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM3_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM3_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM3_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM3_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM3_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM3_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM3_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM3_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM3_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM3_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM3_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM3_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM3_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM3_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM3_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM3_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM3_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM3_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM3_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM3_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM3_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM3_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM3_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM3_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM3_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM3_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM3_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM3_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM3_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM3_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM3_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM3_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM3_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM3_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM3_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM3_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM3_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM3_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM3_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM3_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM3_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM3_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM3_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM3_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM3_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM3_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM3_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM3_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM3_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM3_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM3_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM3_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM3_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM3_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(3), SSR=>'0', WE=>we, DO=>DOvec(3)(15 downto 8), DOP=>open);
RAM3_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM3_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM3_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM3_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM3_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM3_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM3_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM3_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM3_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM3_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM3_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM3_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM3_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM3_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM3_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM3_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM3_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM3_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM3_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM3_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM3_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM3_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM3_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM3_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM3_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM3_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM3_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM3_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM3_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM3_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM3_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM3_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM3_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM3_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM3_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM3_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM3_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM3_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM3_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM3_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM3_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM3_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM3_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM3_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM3_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM3_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM3_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM3_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM3_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM3_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM3_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM3_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM3_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM3_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM3_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM3_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM3_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM3_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM3_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM3_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM3_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM3_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM3_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM3_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM3_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(3), SSR=>'0', WE=>we, DO=>DOvec(3)(23 downto 16), DOP=>open);


RAM4_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM4_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM4_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM4_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM4_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM4_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM4_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM4_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM4_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM4_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM4_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM4_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM4_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM4_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM4_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM4_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM4_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM4_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM4_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM4_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM4_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM4_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM4_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM4_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM4_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM4_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM4_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM4_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM4_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM4_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM4_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM4_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM4_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM4_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM4_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM4_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM4_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM4_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM4_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM4_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM4_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM4_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM4_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM4_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM4_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM4_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM4_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM4_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM4_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM4_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM4_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM4_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM4_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM4_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM4_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM4_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM4_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM4_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM4_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM4_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM4_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM4_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM4_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM4_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM4_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(4), SSR=>'0', WE=>we, DO=>DOvec(4)(7 downto 0), DOP=>open);
RAM4_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM4_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM4_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM4_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM4_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM4_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM4_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM4_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM4_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM4_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM4_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM4_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM4_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM4_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM4_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM4_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM4_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM4_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM4_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM4_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM4_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM4_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM4_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM4_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM4_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM4_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM4_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM4_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM4_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM4_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM4_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM4_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM4_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM4_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM4_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM4_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM4_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM4_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM4_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM4_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM4_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM4_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM4_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM4_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM4_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM4_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM4_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM4_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM4_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM4_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM4_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM4_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM4_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM4_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM4_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM4_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM4_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM4_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM4_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM4_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM4_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM4_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM4_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM4_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM4_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(4), SSR=>'0', WE=>we, DO=>DOvec(4)(15 downto 8), DOP=>open);
RAM4_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM4_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM4_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM4_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM4_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM4_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM4_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM4_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM4_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM4_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM4_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM4_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM4_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM4_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM4_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM4_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM4_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM4_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM4_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM4_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM4_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM4_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM4_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM4_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM4_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM4_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM4_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM4_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM4_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM4_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM4_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM4_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM4_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM4_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM4_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM4_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM4_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM4_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM4_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM4_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM4_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM4_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM4_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM4_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM4_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM4_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM4_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM4_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM4_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM4_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM4_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM4_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM4_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM4_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM4_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM4_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM4_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM4_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM4_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM4_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM4_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM4_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM4_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM4_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM4_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(4), SSR=>'0', WE=>we, DO=>DOvec(4)(23 downto 16), DOP=>open);


RAM5_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM5_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM5_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM5_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM5_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM5_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM5_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM5_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM5_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM5_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM5_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM5_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM5_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM5_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM5_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM5_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM5_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM5_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM5_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM5_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM5_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM5_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM5_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM5_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM5_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM5_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM5_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM5_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM5_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM5_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM5_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM5_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM5_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM5_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM5_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM5_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM5_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM5_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM5_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM5_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM5_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM5_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM5_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM5_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM5_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM5_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM5_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM5_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM5_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM5_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM5_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM5_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM5_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM5_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM5_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM5_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM5_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM5_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM5_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM5_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM5_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM5_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM5_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM5_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM5_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(5), SSR=>'0', WE=>we, DO=>DOvec(5)(7 downto 0), DOP=>open);
RAM5_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM5_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM5_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM5_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM5_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM5_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM5_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM5_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM5_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM5_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM5_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM5_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM5_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM5_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM5_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM5_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM5_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM5_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM5_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM5_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM5_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM5_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM5_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM5_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM5_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM5_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM5_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM5_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM5_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM5_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM5_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM5_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM5_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM5_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM5_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM5_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM5_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM5_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM5_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM5_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM5_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM5_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM5_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM5_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM5_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM5_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM5_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM5_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM5_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM5_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM5_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM5_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM5_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM5_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM5_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM5_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM5_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM5_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM5_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM5_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM5_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM5_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM5_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM5_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM5_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(5), SSR=>'0', WE=>we, DO=>DOvec(5)(15 downto 8), DOP=>open);
RAM5_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM5_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM5_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM5_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM5_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM5_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM5_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM5_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM5_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM5_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM5_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM5_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM5_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM5_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM5_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM5_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM5_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM5_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM5_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM5_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM5_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM5_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM5_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM5_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM5_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM5_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM5_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM5_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM5_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM5_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM5_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM5_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM5_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM5_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM5_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM5_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM5_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM5_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM5_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM5_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM5_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM5_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM5_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM5_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM5_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM5_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM5_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM5_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM5_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM5_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM5_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM5_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM5_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM5_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM5_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM5_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM5_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM5_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM5_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM5_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM5_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM5_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM5_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM5_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM5_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(5), SSR=>'0', WE=>we, DO=>DOvec(5)(23 downto 16), DOP=>open);


RAM6_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM6_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM6_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM6_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM6_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM6_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM6_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM6_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM6_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM6_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM6_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM6_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM6_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM6_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM6_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM6_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM6_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM6_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM6_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM6_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM6_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM6_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM6_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM6_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM6_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM6_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM6_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM6_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM6_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM6_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM6_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM6_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM6_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM6_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM6_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM6_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM6_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM6_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM6_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM6_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM6_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM6_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM6_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM6_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM6_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM6_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM6_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM6_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM6_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM6_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM6_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM6_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM6_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM6_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM6_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM6_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM6_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM6_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM6_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM6_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM6_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM6_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM6_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM6_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM6_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(6), SSR=>'0', WE=>we, DO=>DOvec(6)(7 downto 0), DOP=>open);
RAM6_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM6_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM6_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM6_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM6_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM6_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM6_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM6_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM6_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM6_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM6_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM6_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM6_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM6_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM6_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM6_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM6_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM6_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM6_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM6_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM6_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM6_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM6_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM6_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM6_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM6_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM6_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM6_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM6_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM6_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM6_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM6_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM6_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM6_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM6_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM6_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM6_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM6_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM6_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM6_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM6_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM6_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM6_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM6_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM6_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM6_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM6_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM6_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM6_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM6_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM6_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM6_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM6_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM6_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM6_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM6_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM6_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM6_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM6_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM6_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM6_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM6_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM6_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM6_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM6_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(6), SSR=>'0', WE=>we, DO=>DOvec(6)(15 downto 8), DOP=>open);
RAM6_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM6_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM6_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM6_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM6_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM6_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM6_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM6_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM6_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM6_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM6_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM6_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM6_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM6_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM6_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM6_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM6_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM6_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM6_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM6_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM6_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM6_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM6_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM6_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM6_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM6_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM6_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM6_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM6_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM6_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM6_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM6_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM6_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM6_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM6_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM6_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM6_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM6_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM6_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM6_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM6_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM6_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM6_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM6_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM6_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM6_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM6_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM6_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM6_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM6_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM6_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM6_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM6_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM6_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM6_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM6_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM6_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM6_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM6_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM6_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM6_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM6_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM6_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM6_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM6_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(6), SSR=>'0', WE=>we, DO=>DOvec(6)(23 downto 16), DOP=>open);


RAM7_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM7_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM7_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM7_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM7_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM7_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM7_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM7_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM7_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM7_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM7_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM7_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM7_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM7_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM7_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM7_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM7_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM7_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM7_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM7_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM7_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM7_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM7_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM7_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM7_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM7_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM7_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM7_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM7_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM7_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM7_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM7_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM7_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM7_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM7_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM7_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM7_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM7_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM7_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM7_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM7_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM7_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM7_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM7_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM7_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM7_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM7_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM7_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM7_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM7_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM7_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM7_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM7_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM7_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM7_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM7_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM7_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM7_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM7_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM7_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM7_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM7_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM7_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM7_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM7_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(7), SSR=>'0', WE=>we, DO=>DOvec(7)(7 downto 0), DOP=>open);
RAM7_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM7_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM7_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM7_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM7_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM7_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM7_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM7_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM7_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM7_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM7_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM7_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM7_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM7_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM7_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM7_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM7_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM7_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM7_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM7_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM7_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM7_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM7_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM7_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM7_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM7_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM7_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM7_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM7_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM7_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM7_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM7_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM7_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM7_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM7_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM7_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM7_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM7_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM7_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM7_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM7_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM7_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM7_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM7_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM7_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM7_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM7_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM7_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM7_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM7_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM7_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM7_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM7_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM7_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM7_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM7_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM7_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM7_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM7_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM7_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM7_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM7_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM7_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM7_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM7_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(7), SSR=>'0', WE=>we, DO=>DOvec(7)(15 downto 8), DOP=>open);
RAM7_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM7_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM7_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM7_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM7_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM7_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM7_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM7_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM7_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM7_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM7_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM7_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM7_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM7_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM7_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM7_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM7_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM7_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM7_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM7_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM7_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM7_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM7_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM7_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM7_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM7_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM7_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM7_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM7_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM7_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM7_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM7_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM7_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM7_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM7_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM7_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM7_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM7_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM7_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM7_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM7_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM7_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM7_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM7_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM7_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM7_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM7_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM7_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM7_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM7_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM7_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM7_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM7_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM7_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM7_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM7_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM7_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM7_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM7_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM7_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM7_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM7_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM7_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM7_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM7_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(7), SSR=>'0', WE=>we, DO=>DOvec(7)(23 downto 16), DOP=>open);


RAM8_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM8_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM8_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM8_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM8_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM8_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM8_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM8_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM8_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM8_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM8_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM8_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM8_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM8_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM8_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM8_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM8_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM8_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM8_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM8_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM8_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM8_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM8_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM8_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM8_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM8_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM8_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM8_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM8_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM8_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM8_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM8_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM8_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM8_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM8_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM8_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM8_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM8_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM8_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM8_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM8_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM8_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM8_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM8_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM8_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM8_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM8_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM8_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM8_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM8_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM8_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM8_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM8_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM8_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM8_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM8_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM8_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM8_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM8_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM8_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM8_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM8_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM8_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM8_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM8_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(8), SSR=>'0', WE=>we, DO=>DOvec(8)(7 downto 0), DOP=>open);
RAM8_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM8_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM8_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM8_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM8_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM8_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM8_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM8_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM8_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM8_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM8_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM8_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM8_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM8_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM8_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM8_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM8_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM8_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM8_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM8_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM8_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM8_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM8_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM8_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM8_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM8_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM8_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM8_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM8_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM8_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM8_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM8_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM8_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM8_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM8_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM8_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM8_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM8_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM8_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM8_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM8_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM8_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM8_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM8_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM8_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM8_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM8_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM8_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM8_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM8_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM8_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM8_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM8_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM8_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM8_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM8_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM8_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM8_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM8_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM8_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM8_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM8_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM8_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM8_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM8_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(8), SSR=>'0', WE=>we, DO=>DOvec(8)(15 downto 8), DOP=>open);
RAM8_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM8_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM8_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM8_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM8_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM8_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM8_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM8_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM8_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM8_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM8_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM8_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM8_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM8_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM8_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM8_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM8_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM8_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM8_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM8_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM8_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM8_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM8_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM8_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM8_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM8_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM8_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM8_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM8_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM8_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM8_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM8_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM8_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM8_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM8_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM8_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM8_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM8_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM8_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM8_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM8_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM8_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM8_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM8_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM8_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM8_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM8_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM8_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM8_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM8_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM8_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM8_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM8_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM8_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM8_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM8_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM8_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM8_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM8_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM8_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM8_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM8_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM8_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM8_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM8_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(8), SSR=>'0', WE=>we, DO=>DOvec(8)(23 downto 16), DOP=>open);


RAM9_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM9_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM9_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM9_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM9_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM9_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM9_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM9_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM9_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM9_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM9_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM9_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM9_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM9_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM9_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM9_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM9_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM9_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM9_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM9_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM9_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM9_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM9_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM9_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM9_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM9_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM9_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM9_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM9_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM9_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM9_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM9_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM9_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM9_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM9_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM9_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM9_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM9_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM9_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM9_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM9_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM9_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM9_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM9_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM9_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM9_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM9_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM9_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM9_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM9_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM9_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM9_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM9_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM9_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM9_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM9_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM9_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM9_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM9_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM9_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM9_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM9_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM9_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM9_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM9_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(9), SSR=>'0', WE=>we, DO=>DOvec(9)(7 downto 0), DOP=>open);
RAM9_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM9_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM9_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM9_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM9_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM9_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM9_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM9_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM9_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM9_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM9_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM9_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM9_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM9_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM9_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM9_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM9_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM9_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM9_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM9_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM9_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM9_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM9_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM9_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM9_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM9_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM9_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM9_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM9_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM9_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM9_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM9_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM9_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM9_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM9_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM9_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM9_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM9_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM9_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM9_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM9_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM9_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM9_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM9_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM9_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM9_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM9_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM9_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM9_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM9_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM9_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM9_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM9_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM9_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM9_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM9_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM9_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM9_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM9_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM9_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM9_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM9_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM9_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM9_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM9_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(9), SSR=>'0', WE=>we, DO=>DOvec(9)(15 downto 8), DOP=>open);
RAM9_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM9_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM9_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM9_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM9_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM9_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM9_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM9_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM9_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM9_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM9_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM9_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM9_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM9_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM9_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM9_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM9_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM9_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM9_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM9_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM9_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM9_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM9_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM9_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM9_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM9_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM9_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM9_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM9_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM9_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM9_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM9_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM9_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM9_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM9_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM9_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM9_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM9_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM9_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM9_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM9_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM9_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM9_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM9_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM9_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM9_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM9_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM9_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM9_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM9_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM9_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM9_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM9_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM9_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM9_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM9_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM9_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM9_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM9_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM9_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM9_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM9_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM9_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM9_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM9_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(9), SSR=>'0', WE=>we, DO=>DOvec(9)(23 downto 16), DOP=>open);


RAM10_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM10_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM10_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM10_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM10_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM10_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM10_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM10_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM10_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM10_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM10_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM10_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM10_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM10_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM10_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM10_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM10_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM10_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM10_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM10_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM10_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM10_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM10_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM10_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM10_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM10_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM10_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM10_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM10_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM10_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM10_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM10_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM10_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM10_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM10_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM10_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM10_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM10_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM10_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM10_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM10_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM10_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM10_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM10_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM10_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM10_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM10_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM10_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM10_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM10_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM10_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM10_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM10_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM10_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM10_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM10_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM10_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM10_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM10_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM10_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM10_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM10_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM10_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM10_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM10_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(10), SSR=>'0', WE=>we, DO=>DOvec(10)(7 downto 0), DOP=>open);
RAM10_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM10_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM10_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM10_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM10_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM10_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM10_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM10_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM10_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM10_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM10_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM10_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM10_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM10_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM10_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM10_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM10_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM10_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM10_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM10_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM10_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM10_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM10_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM10_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM10_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM10_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM10_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM10_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM10_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM10_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM10_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM10_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM10_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM10_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM10_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM10_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM10_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM10_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM10_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM10_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM10_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM10_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM10_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM10_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM10_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM10_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM10_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM10_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM10_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM10_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM10_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM10_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM10_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM10_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM10_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM10_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM10_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM10_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM10_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM10_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM10_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM10_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM10_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM10_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM10_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(10), SSR=>'0', WE=>we, DO=>DOvec(10)(15 downto 8), DOP=>open);
RAM10_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM10_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM10_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM10_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM10_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM10_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM10_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM10_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM10_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM10_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM10_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM10_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM10_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM10_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM10_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM10_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM10_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM10_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM10_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM10_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM10_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM10_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM10_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM10_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM10_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM10_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM10_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM10_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM10_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM10_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM10_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM10_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM10_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM10_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM10_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM10_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM10_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM10_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM10_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM10_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM10_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM10_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM10_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM10_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM10_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM10_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM10_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM10_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM10_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM10_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM10_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM10_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM10_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM10_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM10_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM10_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM10_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM10_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM10_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM10_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM10_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM10_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM10_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM10_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM10_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(10), SSR=>'0', WE=>we, DO=>DOvec(10)(23 downto 16), DOP=>open);


RAM11_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM11_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM11_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM11_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM11_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM11_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM11_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM11_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM11_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM11_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM11_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM11_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM11_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM11_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM11_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM11_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM11_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM11_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM11_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM11_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM11_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM11_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM11_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM11_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM11_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM11_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM11_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM11_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM11_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM11_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM11_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM11_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM11_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM11_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM11_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM11_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM11_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM11_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM11_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM11_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM11_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM11_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM11_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM11_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM11_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM11_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM11_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM11_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM11_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM11_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM11_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM11_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM11_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM11_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM11_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM11_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM11_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM11_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM11_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM11_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM11_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM11_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM11_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM11_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM11_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(11), SSR=>'0', WE=>we, DO=>DOvec(11)(7 downto 0), DOP=>open);
RAM11_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM11_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM11_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM11_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM11_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM11_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM11_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM11_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM11_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM11_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM11_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM11_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM11_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM11_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM11_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM11_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM11_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM11_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM11_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM11_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM11_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM11_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM11_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM11_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM11_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM11_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM11_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM11_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM11_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM11_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM11_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM11_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM11_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM11_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM11_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM11_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM11_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM11_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM11_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM11_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM11_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM11_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM11_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM11_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM11_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM11_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM11_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM11_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM11_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM11_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM11_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM11_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM11_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM11_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM11_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM11_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM11_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM11_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM11_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM11_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM11_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM11_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM11_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM11_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM11_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(11), SSR=>'0', WE=>we, DO=>DOvec(11)(15 downto 8), DOP=>open);
RAM11_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM11_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM11_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM11_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM11_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM11_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM11_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM11_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM11_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM11_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM11_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM11_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM11_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM11_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM11_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM11_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM11_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM11_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM11_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM11_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM11_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM11_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM11_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM11_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM11_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM11_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM11_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM11_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM11_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM11_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM11_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM11_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM11_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM11_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM11_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM11_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM11_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM11_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM11_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM11_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM11_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM11_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM11_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM11_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM11_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM11_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM11_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM11_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM11_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM11_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM11_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM11_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM11_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM11_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM11_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM11_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM11_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM11_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM11_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM11_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM11_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM11_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM11_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM11_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM11_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(11), SSR=>'0', WE=>we, DO=>DOvec(11)(23 downto 16), DOP=>open);


RAM12_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM12_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM12_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM12_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM12_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM12_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM12_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM12_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM12_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM12_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM12_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM12_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM12_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM12_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM12_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM12_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM12_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM12_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM12_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM12_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM12_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM12_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM12_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM12_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM12_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM12_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM12_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM12_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM12_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM12_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM12_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM12_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM12_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM12_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM12_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM12_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM12_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM12_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM12_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM12_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM12_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM12_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM12_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM12_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM12_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM12_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM12_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM12_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM12_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM12_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM12_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM12_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM12_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM12_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM12_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM12_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM12_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM12_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM12_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM12_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM12_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM12_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM12_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM12_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM12_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(12), SSR=>'0', WE=>we, DO=>DOvec(12)(7 downto 0), DOP=>open);
RAM12_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM12_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM12_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM12_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM12_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM12_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM12_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM12_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM12_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM12_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM12_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM12_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM12_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM12_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM12_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM12_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM12_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM12_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM12_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM12_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM12_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM12_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM12_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM12_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM12_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM12_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM12_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM12_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM12_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM12_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM12_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM12_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM12_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM12_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM12_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM12_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM12_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM12_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM12_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM12_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM12_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM12_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM12_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM12_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM12_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM12_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM12_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM12_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM12_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM12_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM12_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM12_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM12_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM12_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM12_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM12_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM12_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM12_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM12_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM12_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM12_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM12_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM12_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM12_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM12_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(12), SSR=>'0', WE=>we, DO=>DOvec(12)(15 downto 8), DOP=>open);
RAM12_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM12_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM12_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM12_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM12_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM12_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM12_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM12_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM12_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM12_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM12_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM12_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM12_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM12_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM12_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM12_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM12_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM12_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM12_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM12_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM12_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM12_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM12_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM12_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM12_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM12_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM12_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM12_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM12_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM12_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM12_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM12_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM12_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM12_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM12_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM12_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM12_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM12_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM12_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM12_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM12_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM12_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM12_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM12_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM12_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM12_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM12_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM12_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM12_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM12_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM12_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM12_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM12_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM12_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM12_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM12_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM12_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM12_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM12_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM12_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM12_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM12_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM12_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM12_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM12_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(12), SSR=>'0', WE=>we, DO=>DOvec(12)(23 downto 16), DOP=>open);


RAM13_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM13_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM13_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM13_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM13_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM13_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM13_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM13_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM13_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM13_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM13_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM13_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM13_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM13_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM13_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM13_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM13_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM13_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM13_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM13_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM13_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM13_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM13_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM13_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM13_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM13_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM13_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM13_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM13_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM13_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM13_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM13_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM13_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM13_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM13_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM13_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM13_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM13_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM13_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM13_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM13_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM13_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM13_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM13_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM13_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM13_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM13_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM13_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM13_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM13_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM13_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM13_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM13_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM13_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM13_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM13_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM13_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM13_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM13_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM13_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM13_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM13_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM13_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM13_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM13_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(13), SSR=>'0', WE=>we, DO=>DOvec(13)(7 downto 0), DOP=>open);
RAM13_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM13_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM13_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM13_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM13_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM13_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM13_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM13_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM13_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM13_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM13_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM13_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM13_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM13_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM13_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM13_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM13_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM13_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM13_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM13_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM13_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM13_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM13_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM13_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM13_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM13_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM13_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM13_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM13_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM13_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM13_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM13_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM13_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM13_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM13_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM13_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM13_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM13_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM13_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM13_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM13_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM13_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM13_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM13_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM13_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM13_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM13_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM13_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM13_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM13_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM13_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM13_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM13_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM13_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM13_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM13_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM13_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM13_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM13_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM13_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM13_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM13_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM13_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM13_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM13_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(13), SSR=>'0', WE=>we, DO=>DOvec(13)(15 downto 8), DOP=>open);
RAM13_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM13_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM13_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM13_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM13_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM13_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM13_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM13_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM13_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM13_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM13_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM13_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM13_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM13_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM13_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM13_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM13_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM13_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM13_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM13_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM13_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM13_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM13_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM13_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM13_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM13_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM13_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM13_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM13_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM13_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM13_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM13_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM13_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM13_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM13_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM13_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM13_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM13_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM13_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM13_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM13_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM13_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM13_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM13_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM13_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM13_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM13_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM13_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM13_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM13_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM13_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM13_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM13_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM13_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM13_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM13_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM13_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM13_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM13_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM13_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM13_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM13_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM13_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM13_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM13_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(13), SSR=>'0', WE=>we, DO=>DOvec(13)(23 downto 16), DOP=>open);


RAM14_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM14_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM14_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM14_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM14_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM14_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM14_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM14_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM14_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM14_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM14_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM14_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM14_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM14_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM14_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM14_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM14_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM14_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM14_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM14_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM14_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM14_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM14_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM14_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM14_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM14_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM14_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM14_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM14_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM14_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM14_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM14_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM14_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM14_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM14_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM14_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM14_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM14_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM14_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM14_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM14_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM14_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM14_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM14_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM14_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM14_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM14_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM14_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM14_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM14_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM14_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM14_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM14_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM14_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM14_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM14_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM14_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM14_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM14_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM14_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM14_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM14_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM14_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM14_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM14_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(14), SSR=>'0', WE=>we, DO=>DOvec(14)(7 downto 0), DOP=>open);
RAM14_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM14_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM14_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM14_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM14_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM14_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM14_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM14_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM14_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM14_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM14_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM14_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM14_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM14_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM14_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM14_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM14_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM14_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM14_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM14_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM14_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM14_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM14_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM14_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM14_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM14_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM14_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM14_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM14_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM14_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM14_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM14_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM14_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM14_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM14_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM14_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM14_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM14_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM14_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM14_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM14_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM14_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM14_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM14_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM14_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM14_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM14_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM14_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM14_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM14_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM14_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM14_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM14_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM14_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM14_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM14_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM14_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM14_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM14_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM14_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM14_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM14_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM14_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM14_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM14_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(14), SSR=>'0', WE=>we, DO=>DOvec(14)(15 downto 8), DOP=>open);
RAM14_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM14_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM14_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM14_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM14_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM14_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM14_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM14_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM14_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM14_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM14_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM14_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM14_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM14_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM14_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM14_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM14_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM14_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM14_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM14_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM14_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM14_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM14_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM14_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM14_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM14_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM14_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM14_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM14_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM14_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM14_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM14_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM14_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM14_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM14_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM14_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM14_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM14_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM14_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM14_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM14_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM14_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM14_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM14_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM14_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM14_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM14_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM14_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM14_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM14_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM14_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM14_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM14_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM14_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM14_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM14_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM14_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM14_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM14_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM14_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM14_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM14_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM14_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM14_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM14_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(14), SSR=>'0', WE=>we, DO=>DOvec(14)(23 downto 16), DOP=>open);


RAM15_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM15_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM15_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM15_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM15_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM15_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM15_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM15_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM15_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM15_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM15_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM15_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM15_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM15_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM15_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM15_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM15_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM15_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM15_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM15_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM15_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM15_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM15_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM15_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM15_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM15_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM15_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM15_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM15_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM15_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM15_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM15_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM15_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM15_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM15_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM15_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM15_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM15_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM15_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM15_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM15_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM15_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM15_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM15_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM15_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM15_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM15_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM15_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM15_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM15_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM15_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM15_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM15_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM15_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM15_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM15_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM15_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM15_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM15_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM15_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM15_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM15_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM15_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM15_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM15_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(15), SSR=>'0', WE=>we, DO=>DOvec(15)(7 downto 0), DOP=>open);
RAM15_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM15_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM15_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM15_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM15_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM15_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM15_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM15_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM15_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM15_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM15_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM15_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM15_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM15_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM15_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM15_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM15_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM15_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM15_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM15_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM15_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM15_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM15_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM15_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM15_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM15_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM15_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM15_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM15_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM15_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM15_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM15_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM15_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM15_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM15_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM15_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM15_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM15_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM15_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM15_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM15_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM15_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM15_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM15_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM15_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM15_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM15_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM15_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM15_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM15_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM15_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM15_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM15_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM15_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM15_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM15_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM15_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM15_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM15_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM15_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM15_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM15_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM15_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM15_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM15_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(15), SSR=>'0', WE=>we, DO=>DOvec(15)(15 downto 8), DOP=>open);
RAM15_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM15_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM15_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM15_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM15_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM15_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM15_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM15_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM15_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM15_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM15_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM15_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM15_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM15_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM15_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM15_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM15_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM15_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM15_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM15_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM15_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM15_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM15_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM15_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM15_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM15_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM15_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM15_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM15_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM15_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM15_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM15_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM15_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM15_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM15_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM15_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM15_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM15_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM15_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM15_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM15_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM15_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM15_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM15_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM15_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM15_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM15_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM15_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM15_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM15_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM15_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM15_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM15_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM15_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM15_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM15_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM15_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM15_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM15_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM15_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM15_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM15_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM15_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM15_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM15_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(15), SSR=>'0', WE=>we, DO=>DOvec(15)(23 downto 16), DOP=>open);


RAM16_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM16_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM16_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM16_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM16_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM16_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM16_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM16_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM16_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM16_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM16_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM16_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM16_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM16_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM16_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM16_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM16_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM16_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM16_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM16_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM16_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM16_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM16_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM16_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM16_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM16_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM16_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM16_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM16_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM16_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM16_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM16_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM16_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM16_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM16_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM16_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM16_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM16_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM16_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM16_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM16_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM16_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM16_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM16_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM16_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM16_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM16_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM16_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM16_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM16_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM16_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM16_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM16_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM16_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM16_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM16_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM16_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM16_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM16_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM16_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM16_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM16_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM16_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM16_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM16_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(16), SSR=>'0', WE=>we, DO=>DOvec(16)(7 downto 0), DOP=>open);
RAM16_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM16_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM16_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM16_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM16_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM16_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM16_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM16_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM16_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM16_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM16_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM16_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM16_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM16_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM16_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM16_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM16_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM16_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM16_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM16_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM16_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM16_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM16_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM16_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM16_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM16_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM16_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM16_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM16_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM16_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM16_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM16_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM16_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM16_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM16_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM16_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM16_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM16_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM16_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM16_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM16_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM16_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM16_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM16_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM16_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM16_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM16_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM16_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM16_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM16_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM16_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM16_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM16_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM16_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM16_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM16_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM16_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM16_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM16_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM16_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM16_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM16_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM16_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM16_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM16_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(16), SSR=>'0', WE=>we, DO=>DOvec(16)(15 downto 8), DOP=>open);
RAM16_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM16_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM16_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM16_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM16_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM16_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM16_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM16_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM16_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM16_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM16_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM16_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM16_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM16_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM16_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM16_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM16_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM16_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM16_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM16_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM16_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM16_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM16_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM16_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM16_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM16_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM16_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM16_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM16_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM16_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM16_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM16_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM16_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM16_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM16_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM16_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM16_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM16_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM16_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM16_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM16_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM16_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM16_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM16_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM16_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM16_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM16_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM16_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM16_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM16_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM16_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM16_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM16_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM16_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM16_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM16_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM16_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM16_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM16_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM16_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM16_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM16_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM16_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM16_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM16_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(16), SSR=>'0', WE=>we, DO=>DOvec(16)(23 downto 16), DOP=>open);


RAM17_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM17_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM17_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM17_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM17_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM17_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM17_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM17_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM17_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM17_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM17_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM17_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM17_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM17_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM17_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM17_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM17_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM17_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM17_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM17_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM17_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM17_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM17_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM17_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM17_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM17_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM17_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM17_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM17_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM17_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM17_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM17_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM17_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM17_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM17_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM17_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM17_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM17_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM17_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM17_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM17_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM17_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM17_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM17_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM17_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM17_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM17_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM17_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM17_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM17_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM17_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM17_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM17_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM17_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM17_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM17_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM17_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM17_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM17_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM17_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM17_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM17_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM17_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM17_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM17_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(17), SSR=>'0', WE=>we, DO=>DOvec(17)(7 downto 0), DOP=>open);
RAM17_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM17_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM17_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM17_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM17_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM17_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM17_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM17_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM17_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM17_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM17_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM17_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM17_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM17_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM17_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM17_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM17_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM17_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM17_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM17_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM17_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM17_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM17_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM17_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM17_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM17_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM17_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM17_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM17_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM17_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM17_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM17_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM17_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM17_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM17_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM17_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM17_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM17_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM17_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM17_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM17_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM17_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM17_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM17_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM17_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM17_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM17_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM17_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM17_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM17_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM17_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM17_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM17_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM17_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM17_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM17_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM17_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM17_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM17_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM17_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM17_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM17_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM17_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM17_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM17_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(17), SSR=>'0', WE=>we, DO=>DOvec(17)(15 downto 8), DOP=>open);
RAM17_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM17_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM17_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM17_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM17_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM17_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM17_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM17_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM17_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM17_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM17_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM17_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM17_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM17_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM17_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM17_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM17_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM17_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM17_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM17_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM17_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM17_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM17_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM17_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM17_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM17_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM17_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM17_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM17_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM17_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM17_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM17_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM17_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM17_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM17_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM17_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM17_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM17_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM17_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM17_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM17_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM17_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM17_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM17_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM17_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM17_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM17_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM17_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM17_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM17_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM17_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM17_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM17_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM17_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM17_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM17_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM17_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM17_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM17_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM17_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM17_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM17_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM17_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM17_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM17_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(17), SSR=>'0', WE=>we, DO=>DOvec(17)(23 downto 16), DOP=>open);


RAM18_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM18_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM18_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM18_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM18_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM18_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM18_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM18_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM18_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM18_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM18_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM18_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM18_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM18_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM18_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM18_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM18_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM18_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM18_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM18_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM18_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM18_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM18_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM18_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM18_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM18_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM18_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM18_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM18_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM18_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM18_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM18_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM18_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM18_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM18_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM18_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM18_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM18_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM18_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM18_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM18_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM18_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM18_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM18_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM18_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM18_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM18_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM18_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM18_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM18_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM18_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM18_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM18_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM18_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM18_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM18_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM18_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM18_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM18_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM18_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM18_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM18_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM18_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM18_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM18_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(18), SSR=>'0', WE=>we, DO=>DOvec(18)(7 downto 0), DOP=>open);
RAM18_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM18_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM18_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM18_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM18_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM18_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM18_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM18_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM18_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM18_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM18_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM18_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM18_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM18_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM18_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM18_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM18_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM18_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM18_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM18_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM18_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM18_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM18_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM18_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM18_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM18_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM18_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM18_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM18_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM18_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM18_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM18_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM18_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM18_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM18_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM18_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM18_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM18_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM18_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM18_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM18_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM18_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM18_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM18_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM18_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM18_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM18_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM18_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM18_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM18_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM18_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM18_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM18_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM18_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM18_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM18_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM18_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM18_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM18_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM18_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM18_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM18_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM18_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM18_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM18_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(18), SSR=>'0', WE=>we, DO=>DOvec(18)(15 downto 8), DOP=>open);
RAM18_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM18_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM18_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM18_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM18_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM18_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM18_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM18_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM18_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM18_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM18_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM18_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM18_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM18_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM18_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM18_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM18_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM18_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM18_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM18_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM18_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM18_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM18_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM18_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM18_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM18_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM18_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM18_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM18_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM18_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM18_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM18_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM18_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM18_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM18_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM18_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM18_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM18_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM18_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM18_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM18_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM18_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM18_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM18_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM18_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM18_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM18_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM18_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM18_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM18_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM18_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM18_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM18_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM18_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM18_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM18_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM18_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM18_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM18_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM18_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM18_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM18_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM18_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM18_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM18_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(18), SSR=>'0', WE=>we, DO=>DOvec(18)(23 downto 16), DOP=>open);


RAM19_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM19_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM19_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM19_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM19_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM19_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM19_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM19_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM19_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM19_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM19_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM19_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM19_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM19_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM19_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM19_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM19_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM19_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM19_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM19_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM19_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM19_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM19_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM19_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM19_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM19_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM19_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM19_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM19_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM19_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM19_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM19_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM19_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM19_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM19_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM19_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM19_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM19_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM19_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM19_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM19_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM19_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM19_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM19_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM19_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM19_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM19_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM19_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM19_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM19_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM19_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM19_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM19_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM19_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM19_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM19_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM19_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM19_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM19_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM19_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM19_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM19_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM19_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM19_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM19_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(19), SSR=>'0', WE=>we, DO=>DOvec(19)(7 downto 0), DOP=>open);
RAM19_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM19_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM19_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM19_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM19_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM19_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM19_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM19_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM19_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM19_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM19_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM19_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM19_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM19_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM19_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM19_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM19_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM19_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM19_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM19_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM19_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM19_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM19_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM19_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM19_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM19_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM19_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM19_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM19_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM19_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM19_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM19_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM19_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM19_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM19_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM19_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM19_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM19_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM19_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM19_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM19_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM19_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM19_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM19_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM19_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM19_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM19_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM19_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM19_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM19_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM19_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM19_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM19_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM19_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM19_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM19_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM19_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM19_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM19_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM19_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM19_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM19_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM19_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM19_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM19_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(19), SSR=>'0', WE=>we, DO=>DOvec(19)(15 downto 8), DOP=>open);
RAM19_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM19_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM19_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM19_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM19_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM19_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM19_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM19_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM19_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM19_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM19_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM19_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM19_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM19_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM19_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM19_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM19_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM19_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM19_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM19_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM19_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM19_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM19_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM19_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM19_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM19_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM19_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM19_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM19_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM19_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM19_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM19_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM19_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM19_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM19_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM19_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM19_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM19_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM19_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM19_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM19_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM19_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM19_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM19_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM19_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM19_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM19_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM19_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM19_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM19_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM19_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM19_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM19_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM19_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM19_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM19_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM19_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM19_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM19_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM19_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM19_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM19_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM19_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM19_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM19_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(19), SSR=>'0', WE=>we, DO=>DOvec(19)(23 downto 16), DOP=>open);


RAM20_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM20_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM20_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM20_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM20_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM20_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM20_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM20_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM20_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM20_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM20_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM20_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM20_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM20_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM20_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM20_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM20_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM20_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM20_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM20_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM20_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM20_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM20_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM20_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM20_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM20_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM20_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM20_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM20_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM20_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM20_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM20_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM20_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM20_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM20_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM20_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM20_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM20_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM20_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM20_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM20_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM20_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM20_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM20_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM20_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM20_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM20_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM20_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM20_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM20_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM20_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM20_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM20_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM20_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM20_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM20_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM20_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM20_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM20_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM20_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM20_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM20_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM20_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM20_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM20_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(20), SSR=>'0', WE=>we, DO=>DOvec(20)(7 downto 0), DOP=>open);
RAM20_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM20_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM20_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM20_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM20_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM20_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM20_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM20_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM20_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM20_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM20_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM20_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM20_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM20_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM20_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM20_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM20_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM20_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM20_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM20_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM20_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM20_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM20_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM20_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM20_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM20_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM20_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM20_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM20_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM20_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM20_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM20_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM20_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM20_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM20_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM20_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM20_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM20_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM20_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM20_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM20_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM20_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM20_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM20_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM20_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM20_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM20_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM20_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM20_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM20_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM20_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM20_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM20_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM20_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM20_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM20_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM20_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM20_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM20_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM20_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM20_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM20_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM20_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM20_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM20_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(20), SSR=>'0', WE=>we, DO=>DOvec(20)(15 downto 8), DOP=>open);
RAM20_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM20_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM20_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM20_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM20_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM20_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM20_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM20_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM20_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM20_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM20_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM20_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM20_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM20_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM20_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM20_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM20_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM20_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM20_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM20_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM20_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM20_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM20_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM20_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM20_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM20_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM20_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM20_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM20_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM20_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM20_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM20_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM20_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM20_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM20_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM20_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM20_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM20_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM20_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM20_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM20_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM20_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM20_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM20_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM20_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM20_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM20_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM20_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM20_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM20_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM20_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM20_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM20_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM20_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM20_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM20_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM20_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM20_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM20_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM20_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM20_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM20_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM20_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM20_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM20_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(20), SSR=>'0', WE=>we, DO=>DOvec(20)(23 downto 16), DOP=>open);


RAM21_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM21_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM21_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM21_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM21_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM21_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM21_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM21_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM21_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM21_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM21_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM21_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM21_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM21_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM21_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM21_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM21_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM21_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM21_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM21_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM21_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM21_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM21_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM21_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM21_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM21_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM21_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM21_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM21_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM21_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM21_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM21_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM21_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM21_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM21_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM21_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM21_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM21_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM21_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM21_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM21_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM21_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM21_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM21_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM21_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM21_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM21_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM21_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM21_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM21_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM21_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM21_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM21_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM21_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM21_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM21_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM21_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM21_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM21_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM21_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM21_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM21_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM21_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM21_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM21_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(21), SSR=>'0', WE=>we, DO=>DOvec(21)(7 downto 0), DOP=>open);
RAM21_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM21_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM21_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM21_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM21_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM21_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM21_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM21_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM21_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM21_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM21_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM21_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM21_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM21_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM21_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM21_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM21_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM21_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM21_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM21_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM21_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM21_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM21_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM21_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM21_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM21_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM21_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM21_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM21_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM21_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM21_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM21_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM21_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM21_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM21_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM21_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM21_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM21_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM21_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM21_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM21_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM21_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM21_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM21_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM21_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM21_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM21_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM21_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM21_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM21_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM21_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM21_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM21_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM21_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM21_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM21_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM21_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM21_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM21_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM21_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM21_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM21_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM21_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM21_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM21_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(21), SSR=>'0', WE=>we, DO=>DOvec(21)(15 downto 8), DOP=>open);
RAM21_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM21_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM21_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM21_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM21_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM21_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM21_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM21_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM21_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM21_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM21_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM21_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM21_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM21_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM21_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM21_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM21_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM21_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM21_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM21_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM21_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM21_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM21_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM21_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM21_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM21_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM21_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM21_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM21_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM21_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM21_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM21_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM21_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM21_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM21_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM21_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM21_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM21_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM21_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM21_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM21_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM21_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM21_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM21_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM21_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM21_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM21_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM21_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM21_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM21_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM21_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM21_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM21_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM21_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM21_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM21_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM21_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM21_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM21_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM21_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM21_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM21_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM21_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM21_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM21_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(21), SSR=>'0', WE=>we, DO=>DOvec(21)(23 downto 16), DOP=>open);


RAM22_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM22_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM22_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM22_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM22_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM22_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM22_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM22_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM22_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM22_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM22_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM22_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM22_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM22_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM22_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM22_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM22_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM22_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM22_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM22_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM22_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM22_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM22_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM22_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM22_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM22_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM22_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM22_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM22_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM22_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM22_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM22_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM22_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM22_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM22_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM22_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM22_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM22_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM22_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM22_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM22_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM22_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM22_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM22_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM22_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM22_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM22_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM22_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM22_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM22_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM22_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM22_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM22_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM22_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM22_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM22_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM22_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM22_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM22_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM22_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM22_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM22_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM22_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM22_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM22_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(22), SSR=>'0', WE=>we, DO=>DOvec(22)(7 downto 0), DOP=>open);
RAM22_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM22_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM22_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM22_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM22_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM22_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM22_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM22_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM22_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM22_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM22_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM22_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM22_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM22_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM22_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM22_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM22_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM22_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM22_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM22_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM22_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM22_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM22_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM22_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM22_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM22_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM22_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM22_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM22_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM22_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM22_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM22_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM22_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM22_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM22_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM22_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM22_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM22_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM22_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM22_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM22_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM22_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM22_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM22_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM22_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM22_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM22_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM22_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM22_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM22_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM22_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM22_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM22_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM22_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM22_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM22_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM22_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM22_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM22_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM22_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM22_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM22_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM22_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM22_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM22_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(22), SSR=>'0', WE=>we, DO=>DOvec(22)(15 downto 8), DOP=>open);
RAM22_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM22_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM22_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM22_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM22_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM22_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM22_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM22_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM22_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM22_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM22_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM22_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM22_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM22_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM22_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM22_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM22_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM22_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM22_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM22_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM22_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM22_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM22_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM22_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM22_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM22_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM22_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM22_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM22_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM22_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM22_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM22_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM22_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM22_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM22_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM22_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM22_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM22_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM22_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM22_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM22_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM22_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM22_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM22_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM22_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM22_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM22_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM22_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM22_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM22_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM22_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM22_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM22_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM22_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM22_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM22_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM22_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM22_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM22_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM22_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM22_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM22_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM22_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM22_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM22_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(22), SSR=>'0', WE=>we, DO=>DOvec(22)(23 downto 16), DOP=>open);


RAM23_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM23_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM23_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM23_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM23_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM23_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM23_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM23_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM23_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM23_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM23_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM23_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM23_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM23_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM23_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM23_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM23_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM23_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM23_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM23_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM23_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM23_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM23_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM23_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM23_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM23_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM23_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM23_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM23_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM23_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM23_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM23_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM23_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM23_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM23_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM23_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM23_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM23_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM23_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM23_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM23_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM23_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM23_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM23_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM23_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM23_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM23_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM23_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM23_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM23_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM23_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM23_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM23_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM23_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM23_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM23_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM23_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM23_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM23_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM23_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM23_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM23_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM23_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM23_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM23_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(23), SSR=>'0', WE=>we, DO=>DOvec(23)(7 downto 0), DOP=>open);
RAM23_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM23_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM23_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM23_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM23_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM23_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM23_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM23_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM23_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM23_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM23_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM23_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM23_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM23_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM23_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM23_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM23_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM23_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM23_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM23_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM23_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM23_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM23_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM23_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM23_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM23_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM23_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM23_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM23_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM23_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM23_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM23_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM23_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM23_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM23_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM23_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM23_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM23_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM23_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM23_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM23_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM23_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM23_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM23_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM23_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM23_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM23_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM23_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM23_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM23_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM23_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM23_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM23_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM23_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM23_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM23_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM23_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM23_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM23_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM23_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM23_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM23_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM23_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM23_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM23_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(23), SSR=>'0', WE=>we, DO=>DOvec(23)(15 downto 8), DOP=>open);
RAM23_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM23_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM23_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM23_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM23_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM23_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM23_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM23_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM23_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM23_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM23_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM23_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM23_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM23_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM23_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM23_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM23_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM23_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM23_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM23_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM23_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM23_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM23_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM23_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM23_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM23_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM23_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM23_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM23_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM23_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM23_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM23_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM23_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM23_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM23_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM23_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM23_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM23_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM23_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM23_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM23_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM23_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM23_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM23_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM23_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM23_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM23_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM23_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM23_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM23_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM23_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM23_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM23_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM23_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM23_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM23_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM23_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM23_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM23_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM23_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM23_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM23_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM23_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM23_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM23_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(23), SSR=>'0', WE=>we, DO=>DOvec(23)(23 downto 16), DOP=>open);


RAM24_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM24_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM24_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM24_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM24_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM24_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM24_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM24_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM24_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM24_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM24_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM24_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM24_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM24_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM24_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM24_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM24_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM24_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM24_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM24_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM24_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM24_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM24_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM24_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM24_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM24_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM24_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM24_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM24_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM24_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM24_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM24_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM24_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM24_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM24_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM24_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM24_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM24_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM24_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM24_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM24_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM24_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM24_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM24_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM24_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM24_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM24_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM24_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM24_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM24_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM24_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM24_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM24_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM24_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM24_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM24_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM24_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM24_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM24_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM24_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM24_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM24_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM24_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM24_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM24_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(24), SSR=>'0', WE=>we, DO=>DOvec(24)(7 downto 0), DOP=>open);
RAM24_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM24_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM24_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM24_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM24_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM24_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM24_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM24_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM24_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM24_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM24_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM24_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM24_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM24_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM24_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM24_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM24_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM24_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM24_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM24_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM24_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM24_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM24_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM24_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM24_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM24_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM24_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM24_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM24_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM24_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM24_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM24_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM24_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM24_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM24_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM24_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM24_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM24_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM24_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM24_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM24_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM24_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM24_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM24_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM24_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM24_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM24_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM24_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM24_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM24_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM24_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM24_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM24_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM24_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM24_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM24_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM24_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM24_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM24_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM24_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM24_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM24_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM24_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM24_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM24_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(24), SSR=>'0', WE=>we, DO=>DOvec(24)(15 downto 8), DOP=>open);
RAM24_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM24_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM24_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM24_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM24_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM24_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM24_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM24_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM24_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM24_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM24_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM24_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM24_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM24_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM24_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM24_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM24_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM24_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM24_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM24_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM24_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM24_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM24_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM24_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM24_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM24_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM24_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM24_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM24_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM24_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM24_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM24_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM24_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM24_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM24_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM24_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM24_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM24_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM24_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM24_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM24_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM24_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM24_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM24_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM24_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM24_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM24_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM24_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM24_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM24_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM24_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM24_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM24_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM24_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM24_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM24_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM24_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM24_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM24_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM24_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM24_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM24_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM24_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM24_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM24_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(24), SSR=>'0', WE=>we, DO=>DOvec(24)(23 downto 16), DOP=>open);


RAM25_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM25_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM25_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM25_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM25_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM25_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM25_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM25_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM25_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM25_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM25_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM25_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM25_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM25_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM25_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM25_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM25_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM25_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM25_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM25_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM25_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM25_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM25_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM25_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM25_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM25_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM25_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM25_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM25_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM25_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM25_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM25_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM25_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM25_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM25_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM25_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM25_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM25_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM25_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM25_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM25_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM25_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM25_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM25_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM25_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM25_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM25_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM25_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM25_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM25_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM25_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM25_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM25_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM25_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM25_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM25_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM25_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM25_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM25_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM25_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM25_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM25_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM25_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM25_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM25_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(25), SSR=>'0', WE=>we, DO=>DOvec(25)(7 downto 0), DOP=>open);
RAM25_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM25_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM25_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM25_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM25_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM25_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM25_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM25_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM25_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM25_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM25_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM25_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM25_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM25_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM25_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM25_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM25_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM25_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM25_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM25_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM25_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM25_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM25_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM25_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM25_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM25_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM25_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM25_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM25_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM25_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM25_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM25_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM25_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM25_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM25_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM25_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM25_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM25_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM25_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM25_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM25_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM25_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM25_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM25_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM25_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM25_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM25_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM25_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM25_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM25_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM25_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM25_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM25_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM25_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM25_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM25_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM25_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM25_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM25_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM25_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM25_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM25_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM25_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM25_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM25_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(25), SSR=>'0', WE=>we, DO=>DOvec(25)(15 downto 8), DOP=>open);
RAM25_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM25_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM25_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM25_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM25_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM25_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM25_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM25_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM25_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM25_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM25_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM25_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM25_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM25_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM25_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM25_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM25_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM25_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM25_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM25_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM25_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM25_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM25_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM25_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM25_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM25_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM25_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM25_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM25_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM25_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM25_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM25_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM25_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM25_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM25_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM25_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM25_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM25_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM25_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM25_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM25_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM25_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM25_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM25_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM25_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM25_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM25_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM25_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM25_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM25_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM25_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM25_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM25_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM25_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM25_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM25_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM25_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM25_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM25_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM25_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM25_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM25_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM25_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM25_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM25_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(25), SSR=>'0', WE=>we, DO=>DOvec(25)(23 downto 16), DOP=>open);


RAM26_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM26_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM26_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM26_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM26_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM26_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM26_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM26_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM26_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM26_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM26_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM26_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM26_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM26_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM26_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM26_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM26_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM26_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM26_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM26_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM26_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM26_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM26_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM26_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM26_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM26_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM26_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM26_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM26_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM26_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM26_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM26_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM26_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM26_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM26_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM26_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM26_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM26_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM26_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM26_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM26_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM26_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM26_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM26_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM26_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM26_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM26_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM26_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM26_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM26_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM26_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM26_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM26_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM26_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM26_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM26_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM26_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM26_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM26_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM26_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM26_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM26_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM26_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM26_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM26_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(26), SSR=>'0', WE=>we, DO=>DOvec(26)(7 downto 0), DOP=>open);
RAM26_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM26_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM26_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM26_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM26_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM26_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM26_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM26_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM26_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM26_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM26_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM26_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM26_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM26_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM26_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM26_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM26_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM26_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM26_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM26_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM26_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM26_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM26_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM26_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM26_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM26_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM26_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM26_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM26_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM26_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM26_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM26_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM26_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM26_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM26_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM26_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM26_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM26_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM26_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM26_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM26_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM26_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM26_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM26_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM26_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM26_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM26_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM26_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM26_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM26_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM26_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM26_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM26_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM26_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM26_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM26_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM26_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM26_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM26_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM26_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM26_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM26_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM26_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM26_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM26_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(26), SSR=>'0', WE=>we, DO=>DOvec(26)(15 downto 8), DOP=>open);
RAM26_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM26_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM26_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM26_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM26_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM26_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM26_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM26_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM26_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM26_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM26_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM26_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM26_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM26_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM26_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM26_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM26_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM26_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM26_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM26_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM26_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM26_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM26_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM26_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM26_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM26_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM26_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM26_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM26_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM26_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM26_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM26_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM26_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM26_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM26_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM26_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM26_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM26_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM26_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM26_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM26_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM26_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM26_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM26_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM26_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM26_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM26_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM26_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM26_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM26_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM26_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM26_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM26_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM26_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM26_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM26_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM26_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM26_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM26_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM26_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM26_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM26_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM26_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM26_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM26_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(26), SSR=>'0', WE=>we, DO=>DOvec(26)(23 downto 16), DOP=>open);


RAM27_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM27_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM27_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM27_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM27_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM27_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM27_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM27_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM27_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM27_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM27_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM27_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM27_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM27_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM27_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM27_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM27_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM27_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM27_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM27_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM27_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM27_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM27_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM27_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM27_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM27_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM27_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM27_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM27_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM27_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM27_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM27_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM27_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM27_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM27_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM27_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM27_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM27_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM27_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM27_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM27_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM27_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM27_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM27_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM27_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM27_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM27_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM27_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM27_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM27_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM27_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM27_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM27_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM27_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM27_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM27_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM27_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM27_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM27_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM27_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM27_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM27_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM27_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM27_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM27_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(27), SSR=>'0', WE=>we, DO=>DOvec(27)(7 downto 0), DOP=>open);
RAM27_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM27_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM27_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM27_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM27_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM27_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM27_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM27_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM27_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM27_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM27_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM27_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM27_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM27_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM27_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM27_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM27_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM27_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM27_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM27_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM27_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM27_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM27_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM27_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM27_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM27_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM27_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM27_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM27_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM27_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM27_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM27_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM27_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM27_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM27_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM27_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM27_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM27_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM27_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM27_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM27_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM27_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM27_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM27_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM27_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM27_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM27_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM27_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM27_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM27_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM27_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM27_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM27_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM27_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM27_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM27_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM27_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM27_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM27_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM27_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM27_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM27_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM27_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM27_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM27_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(27), SSR=>'0', WE=>we, DO=>DOvec(27)(15 downto 8), DOP=>open);
RAM27_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM27_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM27_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM27_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM27_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM27_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM27_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM27_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM27_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM27_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM27_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM27_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM27_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM27_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM27_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM27_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM27_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM27_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM27_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM27_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM27_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM27_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM27_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM27_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM27_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM27_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM27_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM27_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM27_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM27_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM27_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM27_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM27_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM27_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM27_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM27_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM27_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM27_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM27_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM27_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM27_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM27_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM27_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM27_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM27_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM27_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM27_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM27_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM27_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM27_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM27_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM27_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM27_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM27_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM27_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM27_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM27_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM27_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM27_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM27_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM27_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM27_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM27_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM27_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM27_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(27), SSR=>'0', WE=>we, DO=>DOvec(27)(23 downto 16), DOP=>open);


RAM28_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM28_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM28_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM28_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM28_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM28_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM28_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM28_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM28_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM28_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM28_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM28_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM28_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM28_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM28_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM28_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM28_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM28_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM28_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM28_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM28_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM28_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM28_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM28_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM28_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM28_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM28_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM28_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM28_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM28_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM28_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM28_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM28_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM28_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM28_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM28_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM28_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM28_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM28_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM28_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM28_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM28_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM28_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM28_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM28_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM28_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM28_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM28_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM28_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM28_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM28_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM28_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM28_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM28_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM28_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM28_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM28_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM28_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM28_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM28_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM28_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM28_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM28_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM28_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM28_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(28), SSR=>'0', WE=>we, DO=>DOvec(28)(7 downto 0), DOP=>open);
RAM28_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM28_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM28_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM28_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM28_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM28_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM28_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM28_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM28_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM28_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM28_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM28_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM28_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM28_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM28_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM28_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM28_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM28_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM28_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM28_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM28_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM28_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM28_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM28_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM28_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM28_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM28_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM28_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM28_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM28_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM28_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM28_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM28_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM28_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM28_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM28_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM28_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM28_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM28_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM28_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM28_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM28_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM28_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM28_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM28_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM28_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM28_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM28_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM28_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM28_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM28_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM28_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM28_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM28_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM28_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM28_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM28_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM28_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM28_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM28_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM28_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM28_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM28_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM28_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM28_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(28), SSR=>'0', WE=>we, DO=>DOvec(28)(15 downto 8), DOP=>open);
RAM28_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM28_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM28_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM28_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM28_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM28_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM28_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM28_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM28_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM28_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM28_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM28_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM28_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM28_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM28_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM28_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM28_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM28_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM28_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM28_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM28_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM28_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM28_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM28_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM28_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM28_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM28_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM28_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM28_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM28_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM28_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM28_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM28_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM28_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM28_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM28_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM28_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM28_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM28_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM28_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM28_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM28_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM28_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM28_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM28_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM28_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM28_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM28_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM28_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM28_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM28_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM28_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM28_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM28_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM28_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM28_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM28_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM28_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM28_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM28_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM28_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM28_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM28_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM28_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM28_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(28), SSR=>'0', WE=>we, DO=>DOvec(28)(23 downto 16), DOP=>open);


RAM29_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM29_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM29_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM29_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM29_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM29_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM29_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM29_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM29_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM29_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM29_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM29_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM29_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM29_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM29_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM29_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM29_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM29_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM29_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM29_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM29_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM29_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM29_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM29_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM29_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM29_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM29_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM29_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM29_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM29_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM29_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM29_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM29_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM29_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM29_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM29_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM29_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM29_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM29_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM29_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM29_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM29_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM29_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM29_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM29_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM29_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM29_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM29_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM29_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM29_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM29_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM29_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM29_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM29_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM29_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM29_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM29_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM29_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM29_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM29_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM29_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM29_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM29_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM29_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM29_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(29), SSR=>'0', WE=>we, DO=>DOvec(29)(7 downto 0), DOP=>open);
RAM29_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM29_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM29_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM29_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM29_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM29_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM29_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM29_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM29_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM29_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM29_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM29_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM29_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM29_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM29_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM29_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM29_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM29_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM29_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM29_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM29_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM29_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM29_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM29_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM29_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM29_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM29_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM29_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM29_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM29_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM29_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM29_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM29_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM29_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM29_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM29_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM29_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM29_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM29_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM29_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM29_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM29_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM29_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM29_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM29_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM29_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM29_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM29_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM29_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM29_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM29_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM29_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM29_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM29_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM29_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM29_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM29_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM29_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM29_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM29_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM29_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM29_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM29_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM29_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM29_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(29), SSR=>'0', WE=>we, DO=>DOvec(29)(15 downto 8), DOP=>open);
RAM29_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM29_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM29_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM29_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM29_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM29_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM29_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM29_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM29_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM29_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM29_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM29_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM29_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM29_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM29_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM29_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM29_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM29_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM29_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM29_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM29_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM29_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM29_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM29_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM29_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM29_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM29_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM29_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM29_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM29_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM29_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM29_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM29_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM29_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM29_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM29_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM29_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM29_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM29_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM29_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM29_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM29_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM29_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM29_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM29_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM29_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM29_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM29_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM29_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM29_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM29_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM29_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM29_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM29_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM29_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM29_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM29_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM29_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM29_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM29_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM29_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM29_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM29_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM29_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM29_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(29), SSR=>'0', WE=>we, DO=>DOvec(29)(23 downto 16), DOP=>open);


RAM30_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM30_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM30_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM30_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM30_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM30_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM30_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM30_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM30_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM30_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM30_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM30_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM30_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM30_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM30_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM30_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM30_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM30_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM30_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM30_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM30_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM30_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM30_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM30_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM30_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM30_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM30_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM30_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM30_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM30_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM30_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM30_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM30_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM30_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM30_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM30_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM30_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM30_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM30_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM30_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM30_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM30_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM30_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM30_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM30_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM30_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM30_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM30_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM30_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM30_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM30_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM30_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM30_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM30_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM30_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM30_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM30_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM30_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM30_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM30_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM30_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM30_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM30_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM30_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM30_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(30), SSR=>'0', WE=>we, DO=>DOvec(30)(7 downto 0), DOP=>open);
RAM30_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM30_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM30_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM30_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM30_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM30_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM30_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM30_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM30_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM30_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM30_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM30_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM30_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM30_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM30_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM30_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM30_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM30_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM30_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM30_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM30_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM30_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM30_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM30_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM30_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM30_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM30_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM30_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM30_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM30_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM30_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM30_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM30_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM30_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM30_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM30_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM30_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM30_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM30_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM30_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM30_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM30_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM30_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM30_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM30_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM30_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM30_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM30_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM30_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM30_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM30_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM30_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM30_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM30_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM30_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM30_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM30_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM30_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM30_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM30_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM30_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM30_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM30_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM30_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM30_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(30), SSR=>'0', WE=>we, DO=>DOvec(30)(15 downto 8), DOP=>open);
RAM30_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM30_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM30_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM30_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM30_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM30_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM30_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM30_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM30_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM30_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM30_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM30_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM30_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM30_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM30_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM30_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM30_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM30_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM30_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM30_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM30_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM30_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM30_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM30_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM30_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM30_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM30_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM30_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM30_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM30_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM30_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM30_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM30_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM30_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM30_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM30_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM30_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM30_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM30_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM30_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM30_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM30_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM30_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM30_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM30_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM30_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM30_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM30_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM30_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM30_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM30_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM30_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM30_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM30_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM30_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM30_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM30_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM30_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM30_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM30_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM30_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM30_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM30_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM30_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM30_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(30), SSR=>'0', WE=>we, DO=>DOvec(30)(23 downto 16), DOP=>open);


RAM31_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM31_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM31_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM31_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM31_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM31_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM31_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM31_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM31_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM31_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM31_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM31_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM31_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM31_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM31_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM31_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM31_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM31_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM31_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM31_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM31_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM31_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM31_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM31_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM31_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM31_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM31_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM31_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM31_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM31_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM31_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM31_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM31_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM31_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM31_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM31_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM31_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM31_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM31_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM31_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM31_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM31_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM31_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM31_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM31_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM31_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM31_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM31_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM31_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM31_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM31_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM31_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM31_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM31_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM31_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM31_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM31_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM31_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM31_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM31_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM31_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM31_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM31_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM31_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM31_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(31), SSR=>'0', WE=>we, DO=>DOvec(31)(7 downto 0), DOP=>open);
RAM31_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM31_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM31_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM31_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM31_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM31_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM31_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM31_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM31_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM31_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM31_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM31_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM31_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM31_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM31_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM31_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM31_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM31_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM31_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM31_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM31_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM31_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM31_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM31_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM31_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM31_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM31_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM31_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM31_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM31_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM31_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM31_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM31_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM31_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM31_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM31_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM31_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM31_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM31_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM31_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM31_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM31_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM31_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM31_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM31_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM31_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM31_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM31_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM31_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM31_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM31_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM31_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM31_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM31_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM31_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM31_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM31_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM31_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM31_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM31_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM31_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM31_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM31_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM31_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM31_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(31), SSR=>'0', WE=>we, DO=>DOvec(31)(15 downto 8), DOP=>open);
RAM31_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM31_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM31_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM31_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM31_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM31_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM31_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM31_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM31_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM31_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM31_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM31_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM31_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM31_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM31_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM31_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM31_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM31_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM31_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM31_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM31_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM31_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM31_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM31_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM31_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM31_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM31_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM31_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM31_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM31_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM31_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM31_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM31_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM31_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM31_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM31_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM31_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM31_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM31_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM31_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM31_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM31_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM31_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM31_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM31_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM31_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM31_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM31_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM31_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM31_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM31_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM31_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM31_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM31_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM31_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM31_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM31_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM31_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM31_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM31_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM31_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM31_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM31_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM31_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM31_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(31), SSR=>'0', WE=>we, DO=>DOvec(31)(23 downto 16), DOP=>open);


RAM32_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM32_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM32_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM32_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM32_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM32_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM32_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM32_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM32_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM32_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM32_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM32_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM32_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM32_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM32_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM32_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM32_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM32_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM32_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM32_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM32_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM32_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM32_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM32_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM32_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM32_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM32_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM32_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM32_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM32_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM32_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM32_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM32_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM32_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM32_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM32_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM32_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM32_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM32_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM32_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM32_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM32_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM32_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM32_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM32_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM32_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM32_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM32_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM32_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM32_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM32_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM32_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM32_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM32_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM32_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM32_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM32_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM32_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM32_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM32_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM32_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM32_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM32_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM32_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM32_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(32), SSR=>'0', WE=>we, DO=>DOvec(32)(7 downto 0), DOP=>open);
RAM32_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM32_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM32_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM32_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM32_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM32_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM32_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM32_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM32_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM32_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM32_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM32_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM32_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM32_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM32_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM32_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM32_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM32_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM32_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM32_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM32_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM32_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM32_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM32_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM32_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM32_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM32_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM32_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM32_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM32_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM32_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM32_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM32_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM32_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM32_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM32_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM32_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM32_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM32_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM32_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM32_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM32_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM32_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM32_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM32_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM32_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM32_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM32_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM32_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM32_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM32_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM32_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM32_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM32_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM32_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM32_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM32_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM32_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM32_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM32_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM32_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM32_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM32_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM32_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM32_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(32), SSR=>'0', WE=>we, DO=>DOvec(32)(15 downto 8), DOP=>open);
RAM32_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM32_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM32_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM32_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM32_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM32_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM32_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM32_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM32_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM32_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM32_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM32_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM32_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM32_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM32_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM32_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM32_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM32_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM32_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM32_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM32_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM32_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM32_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM32_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM32_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM32_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM32_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM32_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM32_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM32_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM32_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM32_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM32_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM32_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM32_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM32_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM32_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM32_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM32_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM32_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM32_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM32_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM32_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM32_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM32_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM32_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM32_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM32_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM32_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM32_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM32_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM32_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM32_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM32_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM32_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM32_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM32_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM32_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM32_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM32_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM32_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM32_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM32_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM32_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM32_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(32), SSR=>'0', WE=>we, DO=>DOvec(32)(23 downto 16), DOP=>open);


RAM33_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM33_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM33_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM33_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM33_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM33_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM33_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM33_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM33_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM33_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM33_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM33_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM33_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM33_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM33_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM33_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM33_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM33_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM33_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM33_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM33_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM33_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM33_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM33_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM33_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM33_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM33_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM33_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM33_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM33_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM33_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM33_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM33_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM33_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM33_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM33_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM33_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM33_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM33_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM33_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM33_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM33_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM33_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM33_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM33_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM33_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM33_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM33_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM33_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM33_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM33_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM33_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM33_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM33_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM33_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM33_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM33_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM33_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM33_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM33_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM33_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM33_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM33_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM33_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM33_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(33), SSR=>'0', WE=>we, DO=>DOvec(33)(7 downto 0), DOP=>open);
RAM33_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM33_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM33_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM33_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM33_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM33_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM33_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM33_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM33_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM33_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM33_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM33_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM33_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM33_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM33_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM33_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM33_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM33_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM33_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM33_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM33_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM33_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM33_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM33_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM33_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM33_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM33_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM33_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM33_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM33_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM33_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM33_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM33_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM33_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM33_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM33_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM33_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM33_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM33_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM33_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM33_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM33_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM33_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM33_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM33_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM33_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM33_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM33_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM33_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM33_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM33_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM33_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM33_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM33_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM33_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM33_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM33_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM33_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM33_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM33_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM33_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM33_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM33_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM33_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM33_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(33), SSR=>'0', WE=>we, DO=>DOvec(33)(15 downto 8), DOP=>open);
RAM33_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM33_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM33_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM33_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM33_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM33_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM33_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM33_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM33_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM33_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM33_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM33_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM33_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM33_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM33_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM33_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM33_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM33_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM33_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM33_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM33_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM33_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM33_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM33_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM33_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM33_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM33_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM33_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM33_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM33_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM33_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM33_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM33_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM33_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM33_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM33_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM33_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM33_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM33_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM33_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM33_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM33_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM33_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM33_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM33_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM33_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM33_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM33_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM33_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM33_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM33_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM33_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM33_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM33_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM33_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM33_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM33_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM33_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM33_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM33_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM33_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM33_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM33_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM33_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM33_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(33), SSR=>'0', WE=>we, DO=>DOvec(33)(23 downto 16), DOP=>open);


RAM34_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM34_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM34_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM34_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM34_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM34_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM34_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM34_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM34_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM34_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM34_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM34_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM34_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM34_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM34_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM34_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM34_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM34_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM34_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM34_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM34_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM34_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM34_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM34_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM34_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM34_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM34_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM34_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM34_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM34_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM34_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM34_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM34_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM34_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM34_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM34_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM34_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM34_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM34_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM34_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM34_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM34_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM34_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM34_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM34_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM34_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM34_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM34_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM34_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM34_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM34_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM34_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM34_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM34_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM34_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM34_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM34_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM34_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM34_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM34_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM34_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM34_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM34_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM34_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM34_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(34), SSR=>'0', WE=>we, DO=>DOvec(34)(7 downto 0), DOP=>open);
RAM34_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM34_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM34_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM34_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM34_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM34_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM34_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM34_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM34_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM34_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM34_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM34_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM34_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM34_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM34_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM34_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM34_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM34_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM34_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM34_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM34_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM34_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM34_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM34_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM34_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM34_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM34_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM34_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM34_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM34_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM34_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM34_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM34_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM34_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM34_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM34_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM34_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM34_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM34_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM34_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM34_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM34_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM34_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM34_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM34_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM34_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM34_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM34_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM34_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM34_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM34_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM34_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM34_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM34_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM34_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM34_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM34_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM34_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM34_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM34_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM34_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM34_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM34_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM34_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM34_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(34), SSR=>'0', WE=>we, DO=>DOvec(34)(15 downto 8), DOP=>open);
RAM34_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM34_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM34_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM34_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM34_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM34_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM34_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM34_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM34_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM34_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM34_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM34_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM34_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM34_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM34_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM34_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM34_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM34_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM34_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM34_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM34_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM34_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM34_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM34_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM34_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM34_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM34_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM34_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM34_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM34_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM34_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM34_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM34_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM34_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM34_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM34_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM34_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM34_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM34_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM34_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM34_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM34_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM34_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM34_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM34_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM34_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM34_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM34_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM34_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM34_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM34_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM34_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM34_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM34_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM34_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM34_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM34_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM34_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM34_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM34_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM34_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM34_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM34_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM34_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM34_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(34), SSR=>'0', WE=>we, DO=>DOvec(34)(23 downto 16), DOP=>open);


RAM35_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM35_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM35_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM35_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM35_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM35_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM35_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM35_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM35_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM35_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM35_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM35_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM35_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM35_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM35_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM35_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM35_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM35_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM35_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM35_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM35_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM35_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM35_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM35_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM35_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM35_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM35_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM35_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM35_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM35_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM35_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM35_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM35_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM35_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM35_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM35_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM35_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM35_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM35_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM35_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM35_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM35_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM35_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM35_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM35_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM35_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM35_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM35_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM35_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM35_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM35_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM35_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM35_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM35_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM35_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM35_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM35_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM35_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM35_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM35_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM35_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM35_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM35_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM35_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM35_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(35), SSR=>'0', WE=>we, DO=>DOvec(35)(7 downto 0), DOP=>open);
RAM35_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM35_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM35_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM35_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM35_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM35_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM35_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM35_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM35_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM35_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM35_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM35_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM35_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM35_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM35_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM35_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM35_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM35_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM35_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM35_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM35_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM35_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM35_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM35_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM35_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM35_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM35_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM35_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM35_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM35_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM35_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM35_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM35_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM35_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM35_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM35_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM35_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM35_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM35_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM35_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM35_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM35_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM35_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM35_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM35_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM35_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM35_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM35_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM35_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM35_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM35_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM35_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM35_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM35_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM35_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM35_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM35_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM35_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM35_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM35_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM35_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM35_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM35_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM35_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM35_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(35), SSR=>'0', WE=>we, DO=>DOvec(35)(15 downto 8), DOP=>open);
RAM35_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM35_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM35_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM35_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM35_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM35_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM35_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM35_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM35_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM35_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM35_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM35_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM35_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM35_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM35_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM35_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM35_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM35_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM35_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM35_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM35_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM35_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM35_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM35_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM35_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM35_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM35_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM35_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM35_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM35_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM35_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM35_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM35_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM35_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM35_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM35_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM35_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM35_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM35_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM35_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM35_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM35_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM35_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM35_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM35_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM35_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM35_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM35_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM35_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM35_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM35_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM35_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM35_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM35_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM35_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM35_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM35_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM35_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM35_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM35_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM35_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM35_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM35_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM35_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM35_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(35), SSR=>'0', WE=>we, DO=>DOvec(35)(23 downto 16), DOP=>open);


RAM36_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM36_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM36_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM36_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM36_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM36_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM36_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM36_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM36_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM36_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM36_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM36_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM36_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM36_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM36_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM36_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM36_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM36_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM36_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM36_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM36_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM36_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM36_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM36_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM36_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM36_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM36_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM36_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM36_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM36_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM36_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM36_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM36_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM36_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM36_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM36_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM36_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM36_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM36_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM36_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM36_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM36_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM36_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM36_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM36_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM36_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM36_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM36_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM36_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM36_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM36_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM36_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM36_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM36_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM36_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM36_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM36_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM36_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM36_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM36_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM36_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM36_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM36_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM36_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM36_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(36), SSR=>'0', WE=>we, DO=>DOvec(36)(7 downto 0), DOP=>open);
RAM36_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM36_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM36_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM36_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM36_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM36_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM36_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM36_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM36_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM36_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM36_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM36_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM36_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM36_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM36_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM36_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM36_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM36_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM36_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM36_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM36_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM36_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM36_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM36_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM36_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM36_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM36_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM36_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM36_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM36_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM36_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM36_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM36_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM36_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM36_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM36_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM36_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM36_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM36_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM36_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM36_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM36_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM36_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM36_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM36_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM36_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM36_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM36_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM36_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM36_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM36_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM36_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM36_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM36_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM36_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM36_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM36_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM36_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM36_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM36_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM36_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM36_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM36_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM36_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM36_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(36), SSR=>'0', WE=>we, DO=>DOvec(36)(15 downto 8), DOP=>open);
RAM36_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM36_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM36_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM36_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM36_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM36_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM36_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM36_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM36_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM36_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM36_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM36_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM36_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM36_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM36_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM36_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM36_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM36_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM36_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM36_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM36_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM36_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM36_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM36_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM36_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM36_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM36_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM36_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM36_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM36_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM36_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM36_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM36_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM36_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM36_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM36_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM36_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM36_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM36_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM36_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM36_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM36_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM36_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM36_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM36_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM36_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM36_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM36_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM36_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM36_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM36_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM36_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM36_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM36_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM36_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM36_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM36_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM36_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM36_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM36_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM36_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM36_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM36_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM36_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM36_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(36), SSR=>'0', WE=>we, DO=>DOvec(36)(23 downto 16), DOP=>open);


RAM37_0 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM37_0_INIT_00, INIT_01=>cRAM_VIDEO_RAM37_0_INIT_01, INIT_02=>cRAM_VIDEO_RAM37_0_INIT_02, INIT_03=>cRAM_VIDEO_RAM37_0_INIT_03,
INIT_04=>cRAM_VIDEO_RAM37_0_INIT_04, INIT_05=>cRAM_VIDEO_RAM37_0_INIT_05, INIT_06=>cRAM_VIDEO_RAM37_0_INIT_06, INIT_07=>cRAM_VIDEO_RAM37_0_INIT_07,
INIT_08=>cRAM_VIDEO_RAM37_0_INIT_08, INIT_09=>cRAM_VIDEO_RAM37_0_INIT_09, INIT_0a=>cRAM_VIDEO_RAM37_0_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM37_0_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM37_0_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM37_0_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM37_0_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM37_0_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM37_0_INIT_10, INIT_11=>cRAM_VIDEO_RAM37_0_INIT_11, INIT_12=>cRAM_VIDEO_RAM37_0_INIT_12, INIT_13=>cRAM_VIDEO_RAM37_0_INIT_13,
INIT_14=>cRAM_VIDEO_RAM37_0_INIT_14, INIT_15=>cRAM_VIDEO_RAM37_0_INIT_15, INIT_16=>cRAM_VIDEO_RAM37_0_INIT_16, INIT_17=>cRAM_VIDEO_RAM37_0_INIT_17,
INIT_18=>cRAM_VIDEO_RAM37_0_INIT_18, INIT_19=>cRAM_VIDEO_RAM37_0_INIT_19, INIT_1a=>cRAM_VIDEO_RAM37_0_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM37_0_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM37_0_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM37_0_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM37_0_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM37_0_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM37_0_INIT_20, INIT_21=>cRAM_VIDEO_RAM37_0_INIT_21, INIT_22=>cRAM_VIDEO_RAM37_0_INIT_22, INIT_23=>cRAM_VIDEO_RAM37_0_INIT_23,
INIT_24=>cRAM_VIDEO_RAM37_0_INIT_24, INIT_25=>cRAM_VIDEO_RAM37_0_INIT_25, INIT_26=>cRAM_VIDEO_RAM37_0_INIT_26, INIT_27=>cRAM_VIDEO_RAM37_0_INIT_27,
INIT_28=>cRAM_VIDEO_RAM37_0_INIT_28, INIT_29=>cRAM_VIDEO_RAM37_0_INIT_29, INIT_2a=>cRAM_VIDEO_RAM37_0_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM37_0_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM37_0_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM37_0_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM37_0_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM37_0_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM37_0_INIT_30, INIT_31=>cRAM_VIDEO_RAM37_0_INIT_31, INIT_32=>cRAM_VIDEO_RAM37_0_INIT_32, INIT_33=>cRAM_VIDEO_RAM37_0_INIT_33,
INIT_34=>cRAM_VIDEO_RAM37_0_INIT_34, INIT_35=>cRAM_VIDEO_RAM37_0_INIT_35, INIT_36=>cRAM_VIDEO_RAM37_0_INIT_36, INIT_37=>cRAM_VIDEO_RAM37_0_INIT_37,
INIT_38=>cRAM_VIDEO_RAM37_0_INIT_38, INIT_39=>cRAM_VIDEO_RAM37_0_INIT_39, INIT_3a=>cRAM_VIDEO_RAM37_0_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM37_0_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM37_0_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM37_0_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM37_0_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM37_0_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(37), SSR=>'0', WE=>we, DO=>DOvec(37)(7 downto 0), DOP=>open);
RAM37_1 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM37_1_INIT_00, INIT_01=>cRAM_VIDEO_RAM37_1_INIT_01, INIT_02=>cRAM_VIDEO_RAM37_1_INIT_02, INIT_03=>cRAM_VIDEO_RAM37_1_INIT_03,
INIT_04=>cRAM_VIDEO_RAM37_1_INIT_04, INIT_05=>cRAM_VIDEO_RAM37_1_INIT_05, INIT_06=>cRAM_VIDEO_RAM37_1_INIT_06, INIT_07=>cRAM_VIDEO_RAM37_1_INIT_07,
INIT_08=>cRAM_VIDEO_RAM37_1_INIT_08, INIT_09=>cRAM_VIDEO_RAM37_1_INIT_09, INIT_0a=>cRAM_VIDEO_RAM37_1_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM37_1_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM37_1_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM37_1_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM37_1_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM37_1_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM37_1_INIT_10, INIT_11=>cRAM_VIDEO_RAM37_1_INIT_11, INIT_12=>cRAM_VIDEO_RAM37_1_INIT_12, INIT_13=>cRAM_VIDEO_RAM37_1_INIT_13,
INIT_14=>cRAM_VIDEO_RAM37_1_INIT_14, INIT_15=>cRAM_VIDEO_RAM37_1_INIT_15, INIT_16=>cRAM_VIDEO_RAM37_1_INIT_16, INIT_17=>cRAM_VIDEO_RAM37_1_INIT_17,
INIT_18=>cRAM_VIDEO_RAM37_1_INIT_18, INIT_19=>cRAM_VIDEO_RAM37_1_INIT_19, INIT_1a=>cRAM_VIDEO_RAM37_1_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM37_1_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM37_1_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM37_1_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM37_1_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM37_1_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM37_1_INIT_20, INIT_21=>cRAM_VIDEO_RAM37_1_INIT_21, INIT_22=>cRAM_VIDEO_RAM37_1_INIT_22, INIT_23=>cRAM_VIDEO_RAM37_1_INIT_23,
INIT_24=>cRAM_VIDEO_RAM37_1_INIT_24, INIT_25=>cRAM_VIDEO_RAM37_1_INIT_25, INIT_26=>cRAM_VIDEO_RAM37_1_INIT_26, INIT_27=>cRAM_VIDEO_RAM37_1_INIT_27,
INIT_28=>cRAM_VIDEO_RAM37_1_INIT_28, INIT_29=>cRAM_VIDEO_RAM37_1_INIT_29, INIT_2a=>cRAM_VIDEO_RAM37_1_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM37_1_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM37_1_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM37_1_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM37_1_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM37_1_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM37_1_INIT_30, INIT_31=>cRAM_VIDEO_RAM37_1_INIT_31, INIT_32=>cRAM_VIDEO_RAM37_1_INIT_32, INIT_33=>cRAM_VIDEO_RAM37_1_INIT_33,
INIT_34=>cRAM_VIDEO_RAM37_1_INIT_34, INIT_35=>cRAM_VIDEO_RAM37_1_INIT_35, INIT_36=>cRAM_VIDEO_RAM37_1_INIT_36, INIT_37=>cRAM_VIDEO_RAM37_1_INIT_37,
INIT_38=>cRAM_VIDEO_RAM37_1_INIT_38, INIT_39=>cRAM_VIDEO_RAM37_1_INIT_39, INIT_3a=>cRAM_VIDEO_RAM37_1_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM37_1_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM37_1_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM37_1_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM37_1_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM37_1_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(37), SSR=>'0', WE=>we, DO=>DOvec(37)(15 downto 8), DOP=>open);
RAM37_2 : RAMB16_S9
generic map (
INIT_00=>cRAM_VIDEO_RAM37_2_INIT_00, INIT_01=>cRAM_VIDEO_RAM37_2_INIT_01, INIT_02=>cRAM_VIDEO_RAM37_2_INIT_02, INIT_03=>cRAM_VIDEO_RAM37_2_INIT_03,
INIT_04=>cRAM_VIDEO_RAM37_2_INIT_04, INIT_05=>cRAM_VIDEO_RAM37_2_INIT_05, INIT_06=>cRAM_VIDEO_RAM37_2_INIT_06, INIT_07=>cRAM_VIDEO_RAM37_2_INIT_07,
INIT_08=>cRAM_VIDEO_RAM37_2_INIT_08, INIT_09=>cRAM_VIDEO_RAM37_2_INIT_09, INIT_0a=>cRAM_VIDEO_RAM37_2_INIT_0A, INIT_0b=>cRAM_VIDEO_RAM37_2_INIT_0B,
INIT_0c=>cRAM_VIDEO_RAM37_2_INIT_0C, INIT_0d=>cRAM_VIDEO_RAM37_2_INIT_0D, INIT_0e=>cRAM_VIDEO_RAM37_2_INIT_0E, INIT_0f=>cRAM_VIDEO_RAM37_2_INIT_0F,
INIT_10=>cRAM_VIDEO_RAM37_2_INIT_10, INIT_11=>cRAM_VIDEO_RAM37_2_INIT_11, INIT_12=>cRAM_VIDEO_RAM37_2_INIT_12, INIT_13=>cRAM_VIDEO_RAM37_2_INIT_13,
INIT_14=>cRAM_VIDEO_RAM37_2_INIT_14, INIT_15=>cRAM_VIDEO_RAM37_2_INIT_15, INIT_16=>cRAM_VIDEO_RAM37_2_INIT_16, INIT_17=>cRAM_VIDEO_RAM37_2_INIT_17,
INIT_18=>cRAM_VIDEO_RAM37_2_INIT_18, INIT_19=>cRAM_VIDEO_RAM37_2_INIT_19, INIT_1a=>cRAM_VIDEO_RAM37_2_INIT_1A, INIT_1b=>cRAM_VIDEO_RAM37_2_INIT_1B,
INIT_1c=>cRAM_VIDEO_RAM37_2_INIT_1C, INIT_1d=>cRAM_VIDEO_RAM37_2_INIT_1D, INIT_1e=>cRAM_VIDEO_RAM37_2_INIT_1E, INIT_1f=>cRAM_VIDEO_RAM37_2_INIT_1F,
INIT_20=>cRAM_VIDEO_RAM37_2_INIT_20, INIT_21=>cRAM_VIDEO_RAM37_2_INIT_21, INIT_22=>cRAM_VIDEO_RAM37_2_INIT_22, INIT_23=>cRAM_VIDEO_RAM37_2_INIT_23,
INIT_24=>cRAM_VIDEO_RAM37_2_INIT_24, INIT_25=>cRAM_VIDEO_RAM37_2_INIT_25, INIT_26=>cRAM_VIDEO_RAM37_2_INIT_26, INIT_27=>cRAM_VIDEO_RAM37_2_INIT_27,
INIT_28=>cRAM_VIDEO_RAM37_2_INIT_28, INIT_29=>cRAM_VIDEO_RAM37_2_INIT_29, INIT_2a=>cRAM_VIDEO_RAM37_2_INIT_2A, INIT_2b=>cRAM_VIDEO_RAM37_2_INIT_2B,
INIT_2c=>cRAM_VIDEO_RAM37_2_INIT_2C, INIT_2d=>cRAM_VIDEO_RAM37_2_INIT_2D, INIT_2e=>cRAM_VIDEO_RAM37_2_INIT_2E, INIT_2f=>cRAM_VIDEO_RAM37_2_INIT_2F,
INIT_30=>cRAM_VIDEO_RAM37_2_INIT_30, INIT_31=>cRAM_VIDEO_RAM37_2_INIT_31, INIT_32=>cRAM_VIDEO_RAM37_2_INIT_32, INIT_33=>cRAM_VIDEO_RAM37_2_INIT_33,
INIT_34=>cRAM_VIDEO_RAM37_2_INIT_34, INIT_35=>cRAM_VIDEO_RAM37_2_INIT_35, INIT_36=>cRAM_VIDEO_RAM37_2_INIT_36, INIT_37=>cRAM_VIDEO_RAM37_2_INIT_37,
INIT_38=>cRAM_VIDEO_RAM37_2_INIT_38, INIT_39=>cRAM_VIDEO_RAM37_2_INIT_39, INIT_3a=>cRAM_VIDEO_RAM37_2_INIT_3A, INIT_3b=>cRAM_VIDEO_RAM37_2_INIT_3B,
INIT_3c=>cRAM_VIDEO_RAM37_2_INIT_3C, INIT_3d=>cRAM_VIDEO_RAM37_2_INIT_3D, INIT_3e=>cRAM_VIDEO_RAM37_2_INIT_3E, INIT_3f=>cRAM_VIDEO_RAM37_2_INIT_3F)
port map (ADDR=>std_logic_vector(addr(10 downto 0)), CLK=> CLK, DI=>x"00", DIP(0)=>'0', EN=>en(37), SSR=>'0', WE=>we, DO=>DOvec(37)(23 downto 16), DOP=>open);


end Behavioral;
