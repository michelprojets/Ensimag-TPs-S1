library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;
library UNISIM;
use UNISIM.Vcomponents.ALL;
use work.RAM_Video_data_pkg.all;

-- pour une image 320x240 sur 16 bits avec un pixel par adresse

entity RAM_Video is
        port ( 
                 clka  : in    std_logic;   
                 addra : in    unsigned (16 downto 0); 
                 doa   : out   unsigned(15 downto 0);
                 dia   : in   unsigned(15 downto 0);
                 cea   : in   std_logic;
                 wea   : in   std_logic;
                 clkb  : in    std_logic;   
                 addrb : in    unsigned (16 downto 0); 
                 dob   : out   unsigned(15 downto 0)
             );
end RAM_Video;

architecture BEHAVIORAL of RAM_Video is
   signal enA,enB : unsigned(74 downto 0);
   subtype mot is std_logic_vector(15 downto 0);
   type vec is array (natural range 0 to 74) of mot;
   signal DOvecA,DOvecB : vec;
begin
        process (addra(16 downto 10),DOvecA)
                variable i : natural;
        begin
                ena <= (others => '0');
                i:=to_integer(addra(16 downto 10));
                ena(i) <= cea;
                DOA <= unsigned(DOvecA(i));
        end process; 

        process (addrb(16 downto 10),DOvecb)
                variable i : integer;
        begin
                enb <= (others => '0');
                i:=to_integer(addrb(16 downto 10));
                enb(i) <= '1';
                DOb <= unsigned(DOvecB(i));
        end process; 


RAM0 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM0_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM0_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM0_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM0_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM0_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM0_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM0_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM0_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM0_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM0_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM0_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM0_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM0_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM0_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM0_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM0_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM0_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM0_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM0_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM0_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM0_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM0_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM0_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM0_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM0_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM0_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM0_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM0_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM0_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM0_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM0_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM0_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM0_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM0_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM0_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM0_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM0_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM0_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM0_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM0_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM0_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM0_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM0_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM0_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM0_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM0_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM0_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM0_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM0_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM0_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM0_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM0_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM0_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM0_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM0_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM0_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM0_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM0_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM0_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM0_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM0_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM0_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM0_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM0_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(0), SSRA=>'0', WEA=>wea , DOA=>DOvecA(0), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(0), SSRb=>'0', WEb=>'0', DOb=>DOvecB(0), DOPb=>open);

RAM1 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM1_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM1_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM1_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM1_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM1_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM1_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM1_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM1_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM1_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM1_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM1_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM1_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM1_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM1_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM1_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM1_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM1_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM1_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM1_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM1_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM1_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM1_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM1_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM1_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM1_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM1_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM1_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM1_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM1_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM1_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM1_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM1_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM1_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM1_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM1_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM1_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM1_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM1_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM1_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM1_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM1_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM1_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM1_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM1_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM1_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM1_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM1_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM1_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM1_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM1_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM1_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM1_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM1_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM1_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM1_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM1_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM1_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM1_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM1_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM1_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM1_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM1_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM1_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM1_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(1), SSRA=>'0', WEA=>wea , DOA=>DOvecA(1), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(1), SSRb=>'0', WEb=>'0', DOb=>DOvecB(1), DOPb=>open);

RAM2 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM2_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM2_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM2_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM2_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM2_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM2_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM2_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM2_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM2_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM2_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM2_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM2_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM2_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM2_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM2_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM2_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM2_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM2_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM2_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM2_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM2_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM2_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM2_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM2_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM2_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM2_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM2_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM2_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM2_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM2_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM2_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM2_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM2_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM2_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM2_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM2_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM2_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM2_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM2_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM2_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM2_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM2_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM2_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM2_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM2_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM2_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM2_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM2_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM2_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM2_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM2_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM2_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM2_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM2_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM2_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM2_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM2_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM2_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM2_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM2_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM2_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM2_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM2_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM2_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(2), SSRA=>'0', WEA=>wea , DOA=>DOvecA(2), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(2), SSRb=>'0', WEb=>'0', DOb=>DOvecB(2), DOPb=>open);

RAM3 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM3_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM3_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM3_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM3_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM3_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM3_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM3_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM3_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM3_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM3_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM3_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM3_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM3_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM3_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM3_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM3_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM3_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM3_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM3_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM3_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM3_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM3_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM3_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM3_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM3_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM3_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM3_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM3_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM3_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM3_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM3_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM3_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM3_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM3_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM3_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM3_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM3_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM3_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM3_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM3_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM3_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM3_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM3_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM3_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM3_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM3_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM3_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM3_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM3_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM3_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM3_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM3_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM3_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM3_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM3_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM3_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM3_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM3_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM3_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM3_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM3_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM3_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM3_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM3_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(3), SSRA=>'0', WEA=>wea , DOA=>DOvecA(3), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(3), SSRb=>'0', WEb=>'0', DOb=>DOvecB(3), DOPb=>open);

RAM4 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM4_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM4_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM4_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM4_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM4_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM4_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM4_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM4_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM4_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM4_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM4_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM4_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM4_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM4_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM4_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM4_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM4_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM4_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM4_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM4_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM4_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM4_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM4_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM4_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM4_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM4_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM4_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM4_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM4_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM4_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM4_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM4_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM4_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM4_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM4_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM4_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM4_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM4_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM4_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM4_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM4_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM4_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM4_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM4_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM4_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM4_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM4_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM4_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM4_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM4_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM4_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM4_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM4_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM4_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM4_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM4_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM4_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM4_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM4_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM4_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM4_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM4_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM4_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM4_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(4), SSRA=>'0', WEA=>wea , DOA=>DOvecA(4), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(4), SSRb=>'0', WEb=>'0', DOb=>DOvecB(4), DOPb=>open);

RAM5 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM5_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM5_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM5_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM5_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM5_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM5_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM5_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM5_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM5_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM5_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM5_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM5_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM5_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM5_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM5_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM5_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM5_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM5_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM5_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM5_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM5_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM5_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM5_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM5_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM5_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM5_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM5_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM5_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM5_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM5_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM5_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM5_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM5_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM5_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM5_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM5_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM5_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM5_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM5_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM5_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM5_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM5_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM5_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM5_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM5_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM5_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM5_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM5_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM5_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM5_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM5_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM5_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM5_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM5_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM5_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM5_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM5_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM5_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM5_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM5_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM5_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM5_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM5_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM5_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(5), SSRA=>'0', WEA=>wea , DOA=>DOvecA(5), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(5), SSRb=>'0', WEb=>'0', DOb=>DOvecB(5), DOPb=>open);

RAM6 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM6_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM6_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM6_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM6_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM6_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM6_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM6_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM6_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM6_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM6_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM6_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM6_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM6_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM6_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM6_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM6_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM6_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM6_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM6_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM6_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM6_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM6_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM6_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM6_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM6_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM6_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM6_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM6_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM6_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM6_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM6_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM6_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM6_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM6_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM6_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM6_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM6_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM6_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM6_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM6_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM6_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM6_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM6_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM6_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM6_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM6_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM6_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM6_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM6_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM6_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM6_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM6_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM6_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM6_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM6_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM6_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM6_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM6_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM6_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM6_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM6_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM6_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM6_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM6_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(6), SSRA=>'0', WEA=>wea , DOA=>DOvecA(6), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(6), SSRb=>'0', WEb=>'0', DOb=>DOvecB(6), DOPb=>open);

RAM7 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM7_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM7_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM7_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM7_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM7_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM7_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM7_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM7_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM7_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM7_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM7_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM7_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM7_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM7_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM7_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM7_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM7_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM7_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM7_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM7_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM7_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM7_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM7_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM7_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM7_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM7_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM7_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM7_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM7_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM7_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM7_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM7_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM7_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM7_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM7_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM7_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM7_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM7_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM7_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM7_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM7_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM7_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM7_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM7_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM7_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM7_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM7_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM7_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM7_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM7_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM7_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM7_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM7_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM7_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM7_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM7_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM7_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM7_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM7_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM7_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM7_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM7_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM7_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM7_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(7), SSRA=>'0', WEA=>wea , DOA=>DOvecA(7), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(7), SSRb=>'0', WEb=>'0', DOb=>DOvecB(7), DOPb=>open);

RAM8 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM8_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM8_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM8_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM8_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM8_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM8_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM8_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM8_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM8_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM8_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM8_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM8_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM8_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM8_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM8_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM8_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM8_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM8_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM8_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM8_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM8_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM8_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM8_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM8_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM8_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM8_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM8_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM8_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM8_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM8_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM8_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM8_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM8_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM8_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM8_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM8_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM8_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM8_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM8_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM8_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM8_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM8_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM8_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM8_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM8_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM8_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM8_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM8_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM8_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM8_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM8_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM8_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM8_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM8_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM8_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM8_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM8_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM8_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM8_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM8_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM8_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM8_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM8_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM8_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(8), SSRA=>'0', WEA=>wea , DOA=>DOvecA(8), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(8), SSRb=>'0', WEb=>'0', DOb=>DOvecB(8), DOPb=>open);

RAM9 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM9_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM9_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM9_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM9_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM9_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM9_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM9_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM9_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM9_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM9_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM9_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM9_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM9_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM9_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM9_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM9_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM9_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM9_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM9_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM9_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM9_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM9_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM9_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM9_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM9_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM9_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM9_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM9_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM9_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM9_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM9_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM9_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM9_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM9_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM9_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM9_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM9_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM9_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM9_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM9_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM9_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM9_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM9_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM9_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM9_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM9_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM9_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM9_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM9_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM9_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM9_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM9_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM9_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM9_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM9_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM9_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM9_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM9_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM9_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM9_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM9_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM9_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM9_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM9_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(9), SSRA=>'0', WEA=>wea , DOA=>DOvecA(9), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(9), SSRb=>'0', WEb=>'0', DOb=>DOvecB(9), DOPb=>open);

RAM10 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM10_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM10_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM10_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM10_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM10_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM10_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM10_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM10_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM10_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM10_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM10_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM10_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM10_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM10_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM10_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM10_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM10_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM10_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM10_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM10_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM10_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM10_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM10_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM10_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM10_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM10_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM10_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM10_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM10_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM10_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM10_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM10_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM10_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM10_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM10_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM10_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM10_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM10_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM10_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM10_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM10_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM10_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM10_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM10_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM10_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM10_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM10_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM10_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM10_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM10_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM10_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM10_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM10_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM10_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM10_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM10_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM10_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM10_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM10_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM10_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM10_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM10_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM10_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM10_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(10), SSRA=>'0', WEA=>wea , DOA=>DOvecA(10), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(10), SSRb=>'0', WEb=>'0', DOb=>DOvecB(10), DOPb=>open);

RAM11 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM11_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM11_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM11_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM11_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM11_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM11_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM11_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM11_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM11_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM11_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM11_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM11_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM11_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM11_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM11_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM11_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM11_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM11_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM11_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM11_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM11_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM11_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM11_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM11_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM11_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM11_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM11_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM11_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM11_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM11_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM11_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM11_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM11_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM11_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM11_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM11_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM11_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM11_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM11_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM11_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM11_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM11_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM11_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM11_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM11_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM11_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM11_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM11_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM11_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM11_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM11_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM11_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM11_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM11_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM11_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM11_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM11_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM11_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM11_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM11_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM11_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM11_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM11_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM11_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(11), SSRA=>'0', WEA=>wea , DOA=>DOvecA(11), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(11), SSRb=>'0', WEb=>'0', DOb=>DOvecB(11), DOPb=>open);

RAM12 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM12_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM12_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM12_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM12_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM12_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM12_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM12_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM12_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM12_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM12_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM12_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM12_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM12_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM12_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM12_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM12_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM12_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM12_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM12_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM12_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM12_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM12_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM12_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM12_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM12_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM12_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM12_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM12_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM12_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM12_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM12_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM12_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM12_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM12_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM12_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM12_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM12_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM12_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM12_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM12_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM12_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM12_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM12_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM12_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM12_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM12_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM12_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM12_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM12_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM12_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM12_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM12_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM12_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM12_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM12_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM12_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM12_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM12_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM12_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM12_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM12_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM12_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM12_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM12_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(12), SSRA=>'0', WEA=>wea , DOA=>DOvecA(12), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(12), SSRb=>'0', WEb=>'0', DOb=>DOvecB(12), DOPb=>open);

RAM13 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM13_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM13_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM13_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM13_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM13_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM13_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM13_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM13_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM13_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM13_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM13_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM13_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM13_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM13_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM13_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM13_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM13_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM13_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM13_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM13_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM13_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM13_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM13_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM13_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM13_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM13_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM13_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM13_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM13_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM13_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM13_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM13_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM13_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM13_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM13_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM13_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM13_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM13_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM13_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM13_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM13_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM13_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM13_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM13_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM13_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM13_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM13_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM13_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM13_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM13_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM13_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM13_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM13_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM13_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM13_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM13_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM13_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM13_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM13_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM13_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM13_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM13_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM13_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM13_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(13), SSRA=>'0', WEA=>wea , DOA=>DOvecA(13), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(13), SSRb=>'0', WEb=>'0', DOb=>DOvecB(13), DOPb=>open);

RAM14 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM14_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM14_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM14_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM14_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM14_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM14_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM14_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM14_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM14_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM14_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM14_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM14_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM14_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM14_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM14_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM14_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM14_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM14_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM14_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM14_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM14_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM14_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM14_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM14_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM14_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM14_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM14_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM14_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM14_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM14_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM14_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM14_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM14_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM14_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM14_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM14_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM14_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM14_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM14_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM14_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM14_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM14_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM14_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM14_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM14_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM14_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM14_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM14_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM14_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM14_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM14_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM14_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM14_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM14_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM14_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM14_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM14_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM14_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM14_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM14_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM14_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM14_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM14_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM14_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(14), SSRA=>'0', WEA=>wea , DOA=>DOvecA(14), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(14), SSRb=>'0', WEb=>'0', DOb=>DOvecB(14), DOPb=>open);

RAM15 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM15_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM15_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM15_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM15_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM15_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM15_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM15_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM15_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM15_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM15_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM15_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM15_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM15_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM15_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM15_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM15_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM15_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM15_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM15_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM15_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM15_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM15_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM15_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM15_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM15_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM15_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM15_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM15_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM15_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM15_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM15_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM15_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM15_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM15_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM15_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM15_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM15_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM15_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM15_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM15_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM15_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM15_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM15_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM15_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM15_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM15_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM15_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM15_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM15_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM15_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM15_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM15_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM15_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM15_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM15_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM15_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM15_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM15_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM15_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM15_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM15_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM15_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM15_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM15_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(15), SSRA=>'0', WEA=>wea , DOA=>DOvecA(15), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(15), SSRb=>'0', WEb=>'0', DOb=>DOvecB(15), DOPb=>open);

RAM16 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM16_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM16_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM16_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM16_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM16_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM16_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM16_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM16_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM16_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM16_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM16_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM16_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM16_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM16_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM16_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM16_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM16_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM16_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM16_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM16_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM16_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM16_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM16_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM16_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM16_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM16_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM16_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM16_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM16_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM16_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM16_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM16_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM16_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM16_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM16_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM16_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM16_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM16_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM16_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM16_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM16_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM16_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM16_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM16_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM16_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM16_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM16_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM16_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM16_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM16_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM16_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM16_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM16_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM16_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM16_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM16_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM16_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM16_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM16_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM16_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM16_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM16_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM16_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM16_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(16), SSRA=>'0', WEA=>wea , DOA=>DOvecA(16), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(16), SSRb=>'0', WEb=>'0', DOb=>DOvecB(16), DOPb=>open);

RAM17 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM17_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM17_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM17_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM17_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM17_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM17_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM17_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM17_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM17_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM17_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM17_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM17_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM17_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM17_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM17_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM17_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM17_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM17_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM17_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM17_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM17_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM17_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM17_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM17_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM17_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM17_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM17_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM17_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM17_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM17_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM17_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM17_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM17_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM17_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM17_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM17_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM17_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM17_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM17_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM17_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM17_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM17_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM17_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM17_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM17_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM17_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM17_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM17_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM17_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM17_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM17_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM17_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM17_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM17_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM17_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM17_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM17_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM17_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM17_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM17_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM17_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM17_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM17_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM17_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(17), SSRA=>'0', WEA=>wea , DOA=>DOvecA(17), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(17), SSRb=>'0', WEb=>'0', DOb=>DOvecB(17), DOPb=>open);

RAM18 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM18_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM18_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM18_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM18_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM18_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM18_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM18_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM18_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM18_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM18_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM18_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM18_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM18_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM18_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM18_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM18_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM18_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM18_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM18_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM18_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM18_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM18_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM18_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM18_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM18_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM18_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM18_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM18_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM18_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM18_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM18_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM18_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM18_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM18_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM18_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM18_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM18_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM18_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM18_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM18_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM18_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM18_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM18_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM18_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM18_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM18_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM18_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM18_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM18_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM18_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM18_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM18_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM18_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM18_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM18_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM18_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM18_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM18_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM18_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM18_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM18_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM18_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM18_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM18_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(18), SSRA=>'0', WEA=>wea , DOA=>DOvecA(18), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(18), SSRb=>'0', WEb=>'0', DOb=>DOvecB(18), DOPb=>open);

RAM19 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM19_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM19_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM19_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM19_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM19_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM19_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM19_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM19_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM19_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM19_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM19_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM19_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM19_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM19_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM19_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM19_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM19_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM19_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM19_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM19_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM19_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM19_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM19_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM19_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM19_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM19_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM19_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM19_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM19_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM19_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM19_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM19_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM19_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM19_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM19_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM19_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM19_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM19_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM19_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM19_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM19_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM19_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM19_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM19_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM19_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM19_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM19_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM19_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM19_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM19_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM19_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM19_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM19_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM19_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM19_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM19_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM19_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM19_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM19_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM19_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM19_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM19_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM19_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM19_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(19), SSRA=>'0', WEA=>wea , DOA=>DOvecA(19), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(19), SSRb=>'0', WEb=>'0', DOb=>DOvecB(19), DOPb=>open);

RAM20 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM20_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM20_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM20_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM20_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM20_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM20_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM20_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM20_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM20_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM20_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM20_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM20_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM20_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM20_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM20_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM20_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM20_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM20_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM20_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM20_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM20_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM20_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM20_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM20_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM20_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM20_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM20_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM20_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM20_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM20_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM20_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM20_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM20_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM20_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM20_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM20_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM20_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM20_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM20_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM20_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM20_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM20_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM20_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM20_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM20_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM20_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM20_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM20_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM20_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM20_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM20_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM20_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM20_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM20_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM20_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM20_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM20_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM20_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM20_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM20_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM20_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM20_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM20_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM20_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(20), SSRA=>'0', WEA=>wea , DOA=>DOvecA(20), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(20), SSRb=>'0', WEb=>'0', DOb=>DOvecB(20), DOPb=>open);

RAM21 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM21_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM21_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM21_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM21_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM21_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM21_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM21_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM21_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM21_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM21_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM21_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM21_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM21_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM21_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM21_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM21_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM21_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM21_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM21_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM21_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM21_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM21_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM21_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM21_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM21_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM21_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM21_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM21_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM21_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM21_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM21_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM21_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM21_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM21_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM21_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM21_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM21_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM21_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM21_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM21_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM21_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM21_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM21_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM21_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM21_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM21_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM21_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM21_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM21_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM21_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM21_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM21_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM21_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM21_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM21_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM21_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM21_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM21_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM21_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM21_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM21_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM21_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM21_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM21_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(21), SSRA=>'0', WEA=>wea , DOA=>DOvecA(21), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(21), SSRb=>'0', WEb=>'0', DOb=>DOvecB(21), DOPb=>open);

RAM22 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM22_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM22_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM22_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM22_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM22_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM22_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM22_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM22_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM22_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM22_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM22_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM22_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM22_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM22_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM22_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM22_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM22_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM22_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM22_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM22_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM22_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM22_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM22_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM22_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM22_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM22_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM22_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM22_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM22_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM22_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM22_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM22_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM22_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM22_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM22_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM22_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM22_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM22_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM22_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM22_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM22_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM22_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM22_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM22_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM22_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM22_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM22_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM22_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM22_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM22_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM22_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM22_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM22_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM22_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM22_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM22_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM22_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM22_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM22_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM22_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM22_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM22_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM22_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM22_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(22), SSRA=>'0', WEA=>wea , DOA=>DOvecA(22), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(22), SSRb=>'0', WEb=>'0', DOb=>DOvecB(22), DOPb=>open);

RAM23 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM23_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM23_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM23_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM23_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM23_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM23_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM23_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM23_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM23_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM23_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM23_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM23_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM23_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM23_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM23_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM23_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM23_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM23_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM23_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM23_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM23_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM23_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM23_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM23_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM23_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM23_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM23_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM23_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM23_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM23_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM23_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM23_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM23_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM23_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM23_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM23_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM23_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM23_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM23_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM23_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM23_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM23_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM23_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM23_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM23_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM23_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM23_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM23_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM23_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM23_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM23_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM23_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM23_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM23_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM23_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM23_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM23_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM23_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM23_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM23_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM23_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM23_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM23_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM23_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(23), SSRA=>'0', WEA=>wea , DOA=>DOvecA(23), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(23), SSRb=>'0', WEb=>'0', DOb=>DOvecB(23), DOPb=>open);

RAM24 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM24_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM24_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM24_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM24_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM24_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM24_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM24_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM24_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM24_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM24_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM24_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM24_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM24_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM24_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM24_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM24_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM24_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM24_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM24_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM24_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM24_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM24_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM24_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM24_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM24_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM24_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM24_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM24_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM24_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM24_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM24_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM24_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM24_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM24_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM24_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM24_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM24_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM24_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM24_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM24_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM24_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM24_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM24_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM24_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM24_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM24_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM24_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM24_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM24_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM24_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM24_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM24_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM24_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM24_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM24_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM24_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM24_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM24_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM24_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM24_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM24_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM24_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM24_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM24_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(24), SSRA=>'0', WEA=>wea , DOA=>DOvecA(24), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(24), SSRb=>'0', WEb=>'0', DOb=>DOvecB(24), DOPb=>open);

RAM25 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM25_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM25_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM25_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM25_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM25_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM25_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM25_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM25_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM25_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM25_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM25_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM25_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM25_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM25_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM25_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM25_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM25_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM25_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM25_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM25_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM25_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM25_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM25_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM25_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM25_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM25_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM25_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM25_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM25_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM25_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM25_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM25_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM25_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM25_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM25_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM25_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM25_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM25_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM25_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM25_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM25_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM25_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM25_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM25_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM25_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM25_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM25_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM25_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM25_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM25_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM25_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM25_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM25_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM25_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM25_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM25_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM25_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM25_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM25_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM25_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM25_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM25_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM25_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM25_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(25), SSRA=>'0', WEA=>wea , DOA=>DOvecA(25), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(25), SSRb=>'0', WEb=>'0', DOb=>DOvecB(25), DOPb=>open);

RAM26 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM26_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM26_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM26_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM26_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM26_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM26_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM26_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM26_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM26_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM26_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM26_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM26_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM26_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM26_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM26_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM26_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM26_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM26_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM26_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM26_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM26_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM26_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM26_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM26_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM26_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM26_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM26_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM26_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM26_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM26_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM26_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM26_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM26_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM26_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM26_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM26_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM26_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM26_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM26_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM26_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM26_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM26_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM26_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM26_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM26_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM26_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM26_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM26_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM26_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM26_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM26_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM26_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM26_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM26_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM26_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM26_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM26_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM26_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM26_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM26_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM26_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM26_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM26_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM26_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(26), SSRA=>'0', WEA=>wea , DOA=>DOvecA(26), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(26), SSRb=>'0', WEb=>'0', DOb=>DOvecB(26), DOPb=>open);

RAM27 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM27_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM27_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM27_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM27_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM27_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM27_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM27_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM27_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM27_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM27_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM27_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM27_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM27_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM27_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM27_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM27_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM27_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM27_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM27_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM27_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM27_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM27_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM27_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM27_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM27_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM27_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM27_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM27_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM27_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM27_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM27_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM27_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM27_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM27_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM27_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM27_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM27_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM27_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM27_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM27_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM27_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM27_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM27_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM27_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM27_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM27_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM27_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM27_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM27_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM27_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM27_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM27_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM27_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM27_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM27_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM27_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM27_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM27_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM27_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM27_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM27_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM27_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM27_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM27_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(27), SSRA=>'0', WEA=>wea , DOA=>DOvecA(27), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(27), SSRb=>'0', WEb=>'0', DOb=>DOvecB(27), DOPb=>open);

RAM28 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM28_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM28_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM28_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM28_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM28_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM28_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM28_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM28_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM28_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM28_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM28_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM28_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM28_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM28_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM28_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM28_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM28_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM28_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM28_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM28_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM28_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM28_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM28_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM28_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM28_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM28_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM28_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM28_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM28_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM28_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM28_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM28_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM28_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM28_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM28_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM28_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM28_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM28_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM28_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM28_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM28_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM28_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM28_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM28_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM28_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM28_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM28_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM28_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM28_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM28_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM28_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM28_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM28_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM28_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM28_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM28_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM28_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM28_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM28_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM28_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM28_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM28_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM28_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM28_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(28), SSRA=>'0', WEA=>wea , DOA=>DOvecA(28), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(28), SSRb=>'0', WEb=>'0', DOb=>DOvecB(28), DOPb=>open);

RAM29 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM29_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM29_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM29_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM29_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM29_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM29_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM29_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM29_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM29_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM29_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM29_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM29_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM29_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM29_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM29_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM29_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM29_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM29_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM29_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM29_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM29_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM29_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM29_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM29_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM29_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM29_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM29_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM29_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM29_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM29_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM29_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM29_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM29_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM29_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM29_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM29_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM29_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM29_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM29_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM29_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM29_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM29_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM29_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM29_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM29_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM29_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM29_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM29_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM29_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM29_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM29_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM29_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM29_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM29_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM29_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM29_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM29_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM29_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM29_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM29_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM29_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM29_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM29_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM29_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(29), SSRA=>'0', WEA=>wea , DOA=>DOvecA(29), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(29), SSRb=>'0', WEb=>'0', DOb=>DOvecB(29), DOPb=>open);

RAM30 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM30_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM30_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM30_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM30_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM30_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM30_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM30_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM30_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM30_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM30_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM30_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM30_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM30_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM30_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM30_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM30_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM30_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM30_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM30_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM30_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM30_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM30_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM30_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM30_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM30_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM30_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM30_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM30_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM30_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM30_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM30_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM30_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM30_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM30_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM30_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM30_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM30_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM30_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM30_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM30_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM30_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM30_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM30_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM30_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM30_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM30_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM30_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM30_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM30_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM30_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM30_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM30_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM30_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM30_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM30_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM30_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM30_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM30_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM30_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM30_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM30_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM30_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM30_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM30_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(30), SSRA=>'0', WEA=>wea , DOA=>DOvecA(30), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(30), SSRb=>'0', WEb=>'0', DOb=>DOvecB(30), DOPb=>open);

RAM31 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM31_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM31_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM31_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM31_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM31_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM31_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM31_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM31_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM31_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM31_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM31_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM31_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM31_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM31_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM31_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM31_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM31_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM31_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM31_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM31_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM31_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM31_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM31_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM31_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM31_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM31_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM31_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM31_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM31_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM31_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM31_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM31_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM31_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM31_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM31_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM31_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM31_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM31_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM31_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM31_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM31_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM31_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM31_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM31_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM31_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM31_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM31_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM31_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM31_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM31_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM31_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM31_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM31_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM31_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM31_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM31_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM31_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM31_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM31_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM31_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM31_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM31_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM31_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM31_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(31), SSRA=>'0', WEA=>wea , DOA=>DOvecA(31), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(31), SSRb=>'0', WEb=>'0', DOb=>DOvecB(31), DOPb=>open);

RAM32 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM32_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM32_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM32_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM32_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM32_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM32_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM32_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM32_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM32_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM32_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM32_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM32_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM32_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM32_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM32_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM32_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM32_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM32_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM32_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM32_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM32_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM32_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM32_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM32_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM32_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM32_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM32_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM32_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM32_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM32_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM32_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM32_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM32_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM32_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM32_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM32_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM32_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM32_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM32_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM32_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM32_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM32_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM32_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM32_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM32_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM32_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM32_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM32_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM32_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM32_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM32_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM32_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM32_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM32_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM32_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM32_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM32_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM32_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM32_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM32_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM32_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM32_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM32_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM32_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(32), SSRA=>'0', WEA=>wea , DOA=>DOvecA(32), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(32), SSRb=>'0', WEb=>'0', DOb=>DOvecB(32), DOPb=>open);

RAM33 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM33_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM33_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM33_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM33_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM33_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM33_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM33_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM33_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM33_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM33_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM33_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM33_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM33_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM33_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM33_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM33_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM33_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM33_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM33_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM33_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM33_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM33_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM33_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM33_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM33_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM33_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM33_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM33_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM33_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM33_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM33_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM33_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM33_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM33_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM33_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM33_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM33_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM33_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM33_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM33_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM33_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM33_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM33_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM33_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM33_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM33_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM33_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM33_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM33_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM33_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM33_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM33_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM33_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM33_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM33_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM33_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM33_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM33_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM33_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM33_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM33_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM33_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM33_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM33_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(33), SSRA=>'0', WEA=>wea , DOA=>DOvecA(33), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(33), SSRb=>'0', WEb=>'0', DOb=>DOvecB(33), DOPb=>open);

RAM34 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM34_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM34_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM34_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM34_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM34_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM34_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM34_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM34_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM34_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM34_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM34_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM34_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM34_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM34_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM34_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM34_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM34_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM34_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM34_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM34_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM34_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM34_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM34_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM34_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM34_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM34_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM34_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM34_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM34_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM34_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM34_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM34_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM34_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM34_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM34_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM34_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM34_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM34_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM34_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM34_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM34_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM34_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM34_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM34_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM34_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM34_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM34_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM34_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM34_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM34_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM34_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM34_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM34_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM34_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM34_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM34_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM34_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM34_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM34_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM34_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM34_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM34_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM34_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM34_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(34), SSRA=>'0', WEA=>wea , DOA=>DOvecA(34), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(34), SSRb=>'0', WEb=>'0', DOb=>DOvecB(34), DOPb=>open);

RAM35 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM35_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM35_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM35_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM35_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM35_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM35_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM35_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM35_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM35_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM35_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM35_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM35_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM35_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM35_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM35_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM35_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM35_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM35_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM35_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM35_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM35_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM35_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM35_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM35_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM35_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM35_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM35_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM35_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM35_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM35_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM35_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM35_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM35_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM35_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM35_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM35_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM35_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM35_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM35_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM35_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM35_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM35_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM35_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM35_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM35_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM35_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM35_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM35_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM35_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM35_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM35_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM35_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM35_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM35_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM35_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM35_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM35_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM35_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM35_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM35_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM35_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM35_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM35_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM35_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(35), SSRA=>'0', WEA=>wea , DOA=>DOvecA(35), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(35), SSRb=>'0', WEb=>'0', DOb=>DOvecB(35), DOPb=>open);

RAM36 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM36_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM36_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM36_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM36_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM36_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM36_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM36_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM36_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM36_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM36_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM36_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM36_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM36_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM36_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM36_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM36_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM36_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM36_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM36_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM36_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM36_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM36_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM36_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM36_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM36_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM36_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM36_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM36_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM36_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM36_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM36_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM36_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM36_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM36_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM36_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM36_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM36_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM36_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM36_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM36_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM36_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM36_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM36_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM36_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM36_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM36_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM36_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM36_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM36_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM36_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM36_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM36_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM36_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM36_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM36_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM36_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM36_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM36_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM36_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM36_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM36_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM36_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM36_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM36_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(36), SSRA=>'0', WEA=>wea , DOA=>DOvecA(36), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(36), SSRb=>'0', WEb=>'0', DOb=>DOvecB(36), DOPb=>open);

RAM37 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM37_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM37_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM37_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM37_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM37_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM37_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM37_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM37_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM37_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM37_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM37_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM37_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM37_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM37_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM37_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM37_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM37_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM37_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM37_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM37_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM37_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM37_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM37_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM37_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM37_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM37_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM37_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM37_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM37_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM37_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM37_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM37_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM37_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM37_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM37_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM37_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM37_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM37_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM37_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM37_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM37_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM37_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM37_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM37_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM37_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM37_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM37_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM37_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM37_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM37_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM37_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM37_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM37_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM37_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM37_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM37_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM37_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM37_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM37_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM37_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM37_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM37_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM37_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM37_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(37), SSRA=>'0', WEA=>wea , DOA=>DOvecA(37), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(37), SSRb=>'0', WEb=>'0', DOb=>DOvecB(37), DOPb=>open);

RAM38 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM38_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM38_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM38_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM38_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM38_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM38_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM38_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM38_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM38_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM38_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM38_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM38_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM38_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM38_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM38_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM38_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM38_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM38_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM38_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM38_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM38_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM38_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM38_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM38_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM38_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM38_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM38_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM38_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM38_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM38_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM38_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM38_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM38_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM38_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM38_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM38_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM38_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM38_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM38_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM38_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM38_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM38_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM38_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM38_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM38_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM38_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM38_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM38_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM38_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM38_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM38_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM38_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM38_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM38_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM38_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM38_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM38_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM38_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM38_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM38_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM38_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM38_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM38_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM38_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(38), SSRA=>'0', WEA=>wea , DOA=>DOvecA(38), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(38), SSRb=>'0', WEb=>'0', DOb=>DOvecB(38), DOPb=>open);

RAM39 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM39_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM39_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM39_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM39_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM39_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM39_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM39_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM39_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM39_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM39_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM39_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM39_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM39_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM39_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM39_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM39_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM39_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM39_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM39_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM39_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM39_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM39_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM39_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM39_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM39_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM39_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM39_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM39_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM39_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM39_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM39_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM39_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM39_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM39_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM39_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM39_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM39_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM39_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM39_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM39_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM39_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM39_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM39_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM39_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM39_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM39_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM39_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM39_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM39_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM39_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM39_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM39_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM39_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM39_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM39_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM39_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM39_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM39_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM39_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM39_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM39_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM39_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM39_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM39_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(39), SSRA=>'0', WEA=>wea , DOA=>DOvecA(39), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(39), SSRb=>'0', WEb=>'0', DOb=>DOvecB(39), DOPb=>open);

RAM40 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM40_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM40_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM40_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM40_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM40_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM40_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM40_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM40_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM40_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM40_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM40_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM40_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM40_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM40_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM40_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM40_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM40_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM40_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM40_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM40_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM40_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM40_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM40_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM40_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM40_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM40_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM40_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM40_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM40_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM40_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM40_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM40_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM40_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM40_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM40_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM40_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM40_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM40_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM40_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM40_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM40_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM40_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM40_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM40_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM40_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM40_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM40_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM40_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM40_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM40_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM40_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM40_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM40_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM40_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM40_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM40_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM40_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM40_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM40_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM40_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM40_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM40_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM40_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM40_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(40), SSRA=>'0', WEA=>wea , DOA=>DOvecA(40), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(40), SSRb=>'0', WEb=>'0', DOb=>DOvecB(40), DOPb=>open);

RAM41 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM41_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM41_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM41_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM41_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM41_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM41_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM41_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM41_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM41_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM41_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM41_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM41_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM41_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM41_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM41_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM41_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM41_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM41_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM41_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM41_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM41_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM41_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM41_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM41_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM41_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM41_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM41_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM41_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM41_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM41_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM41_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM41_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM41_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM41_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM41_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM41_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM41_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM41_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM41_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM41_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM41_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM41_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM41_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM41_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM41_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM41_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM41_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM41_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM41_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM41_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM41_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM41_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM41_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM41_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM41_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM41_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM41_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM41_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM41_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM41_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM41_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM41_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM41_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM41_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(41), SSRA=>'0', WEA=>wea , DOA=>DOvecA(41), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(41), SSRb=>'0', WEb=>'0', DOb=>DOvecB(41), DOPb=>open);

RAM42 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM42_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM42_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM42_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM42_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM42_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM42_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM42_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM42_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM42_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM42_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM42_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM42_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM42_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM42_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM42_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM42_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM42_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM42_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM42_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM42_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM42_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM42_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM42_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM42_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM42_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM42_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM42_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM42_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM42_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM42_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM42_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM42_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM42_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM42_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM42_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM42_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM42_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM42_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM42_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM42_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM42_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM42_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM42_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM42_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM42_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM42_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM42_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM42_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM42_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM42_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM42_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM42_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM42_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM42_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM42_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM42_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM42_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM42_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM42_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM42_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM42_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM42_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM42_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM42_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(42), SSRA=>'0', WEA=>wea , DOA=>DOvecA(42), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(42), SSRb=>'0', WEb=>'0', DOb=>DOvecB(42), DOPb=>open);

RAM43 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM43_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM43_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM43_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM43_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM43_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM43_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM43_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM43_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM43_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM43_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM43_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM43_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM43_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM43_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM43_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM43_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM43_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM43_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM43_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM43_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM43_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM43_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM43_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM43_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM43_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM43_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM43_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM43_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM43_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM43_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM43_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM43_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM43_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM43_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM43_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM43_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM43_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM43_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM43_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM43_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM43_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM43_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM43_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM43_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM43_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM43_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM43_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM43_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM43_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM43_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM43_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM43_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM43_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM43_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM43_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM43_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM43_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM43_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM43_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM43_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM43_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM43_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM43_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM43_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(43), SSRA=>'0', WEA=>wea , DOA=>DOvecA(43), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(43), SSRb=>'0', WEb=>'0', DOb=>DOvecB(43), DOPb=>open);

RAM44 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM44_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM44_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM44_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM44_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM44_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM44_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM44_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM44_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM44_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM44_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM44_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM44_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM44_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM44_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM44_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM44_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM44_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM44_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM44_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM44_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM44_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM44_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM44_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM44_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM44_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM44_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM44_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM44_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM44_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM44_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM44_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM44_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM44_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM44_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM44_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM44_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM44_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM44_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM44_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM44_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM44_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM44_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM44_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM44_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM44_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM44_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM44_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM44_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM44_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM44_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM44_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM44_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM44_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM44_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM44_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM44_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM44_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM44_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM44_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM44_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM44_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM44_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM44_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM44_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(44), SSRA=>'0', WEA=>wea , DOA=>DOvecA(44), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(44), SSRb=>'0', WEb=>'0', DOb=>DOvecB(44), DOPb=>open);

RAM45 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM45_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM45_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM45_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM45_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM45_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM45_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM45_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM45_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM45_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM45_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM45_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM45_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM45_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM45_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM45_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM45_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM45_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM45_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM45_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM45_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM45_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM45_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM45_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM45_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM45_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM45_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM45_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM45_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM45_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM45_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM45_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM45_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM45_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM45_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM45_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM45_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM45_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM45_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM45_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM45_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM45_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM45_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM45_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM45_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM45_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM45_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM45_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM45_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM45_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM45_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM45_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM45_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM45_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM45_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM45_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM45_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM45_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM45_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM45_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM45_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM45_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM45_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM45_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM45_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(45), SSRA=>'0', WEA=>wea , DOA=>DOvecA(45), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(45), SSRb=>'0', WEb=>'0', DOb=>DOvecB(45), DOPb=>open);

RAM46 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM46_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM46_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM46_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM46_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM46_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM46_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM46_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM46_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM46_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM46_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM46_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM46_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM46_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM46_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM46_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM46_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM46_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM46_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM46_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM46_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM46_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM46_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM46_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM46_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM46_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM46_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM46_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM46_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM46_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM46_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM46_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM46_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM46_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM46_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM46_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM46_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM46_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM46_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM46_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM46_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM46_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM46_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM46_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM46_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM46_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM46_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM46_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM46_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM46_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM46_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM46_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM46_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM46_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM46_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM46_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM46_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM46_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM46_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM46_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM46_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM46_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM46_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM46_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM46_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(46), SSRA=>'0', WEA=>wea , DOA=>DOvecA(46), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(46), SSRb=>'0', WEb=>'0', DOb=>DOvecB(46), DOPb=>open);

RAM47 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM47_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM47_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM47_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM47_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM47_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM47_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM47_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM47_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM47_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM47_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM47_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM47_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM47_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM47_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM47_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM47_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM47_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM47_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM47_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM47_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM47_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM47_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM47_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM47_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM47_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM47_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM47_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM47_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM47_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM47_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM47_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM47_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM47_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM47_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM47_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM47_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM47_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM47_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM47_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM47_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM47_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM47_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM47_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM47_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM47_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM47_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM47_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM47_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM47_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM47_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM47_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM47_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM47_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM47_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM47_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM47_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM47_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM47_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM47_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM47_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM47_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM47_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM47_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM47_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(47), SSRA=>'0', WEA=>wea , DOA=>DOvecA(47), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(47), SSRb=>'0', WEb=>'0', DOb=>DOvecB(47), DOPb=>open);

RAM48 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM48_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM48_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM48_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM48_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM48_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM48_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM48_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM48_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM48_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM48_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM48_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM48_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM48_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM48_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM48_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM48_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM48_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM48_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM48_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM48_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM48_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM48_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM48_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM48_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM48_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM48_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM48_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM48_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM48_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM48_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM48_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM48_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM48_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM48_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM48_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM48_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM48_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM48_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM48_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM48_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM48_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM48_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM48_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM48_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM48_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM48_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM48_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM48_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM48_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM48_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM48_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM48_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM48_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM48_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM48_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM48_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM48_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM48_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM48_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM48_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM48_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM48_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM48_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM48_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(48), SSRA=>'0', WEA=>wea , DOA=>DOvecA(48), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(48), SSRb=>'0', WEb=>'0', DOb=>DOvecB(48), DOPb=>open);

RAM49 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM49_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM49_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM49_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM49_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM49_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM49_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM49_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM49_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM49_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM49_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM49_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM49_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM49_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM49_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM49_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM49_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM49_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM49_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM49_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM49_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM49_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM49_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM49_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM49_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM49_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM49_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM49_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM49_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM49_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM49_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM49_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM49_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM49_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM49_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM49_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM49_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM49_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM49_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM49_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM49_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM49_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM49_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM49_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM49_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM49_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM49_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM49_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM49_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM49_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM49_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM49_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM49_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM49_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM49_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM49_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM49_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM49_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM49_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM49_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM49_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM49_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM49_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM49_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM49_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(49), SSRA=>'0', WEA=>wea , DOA=>DOvecA(49), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(49), SSRb=>'0', WEb=>'0', DOb=>DOvecB(49), DOPb=>open);

RAM50 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM50_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM50_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM50_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM50_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM50_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM50_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM50_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM50_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM50_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM50_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM50_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM50_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM50_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM50_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM50_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM50_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM50_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM50_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM50_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM50_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM50_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM50_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM50_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM50_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM50_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM50_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM50_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM50_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM50_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM50_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM50_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM50_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM50_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM50_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM50_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM50_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM50_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM50_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM50_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM50_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM50_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM50_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM50_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM50_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM50_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM50_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM50_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM50_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM50_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM50_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM50_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM50_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM50_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM50_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM50_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM50_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM50_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM50_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM50_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM50_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM50_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM50_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM50_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM50_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(50), SSRA=>'0', WEA=>wea , DOA=>DOvecA(50), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(50), SSRb=>'0', WEb=>'0', DOb=>DOvecB(50), DOPb=>open);

RAM51 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM51_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM51_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM51_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM51_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM51_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM51_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM51_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM51_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM51_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM51_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM51_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM51_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM51_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM51_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM51_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM51_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM51_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM51_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM51_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM51_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM51_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM51_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM51_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM51_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM51_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM51_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM51_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM51_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM51_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM51_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM51_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM51_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM51_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM51_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM51_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM51_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM51_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM51_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM51_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM51_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM51_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM51_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM51_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM51_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM51_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM51_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM51_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM51_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM51_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM51_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM51_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM51_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM51_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM51_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM51_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM51_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM51_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM51_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM51_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM51_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM51_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM51_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM51_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM51_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(51), SSRA=>'0', WEA=>wea , DOA=>DOvecA(51), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(51), SSRb=>'0', WEb=>'0', DOb=>DOvecB(51), DOPb=>open);

RAM52 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM52_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM52_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM52_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM52_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM52_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM52_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM52_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM52_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM52_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM52_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM52_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM52_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM52_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM52_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM52_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM52_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM52_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM52_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM52_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM52_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM52_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM52_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM52_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM52_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM52_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM52_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM52_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM52_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM52_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM52_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM52_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM52_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM52_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM52_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM52_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM52_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM52_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM52_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM52_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM52_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM52_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM52_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM52_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM52_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM52_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM52_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM52_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM52_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM52_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM52_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM52_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM52_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM52_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM52_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM52_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM52_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM52_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM52_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM52_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM52_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM52_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM52_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM52_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM52_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(52), SSRA=>'0', WEA=>wea , DOA=>DOvecA(52), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(52), SSRb=>'0', WEb=>'0', DOb=>DOvecB(52), DOPb=>open);

RAM53 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM53_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM53_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM53_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM53_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM53_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM53_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM53_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM53_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM53_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM53_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM53_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM53_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM53_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM53_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM53_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM53_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM53_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM53_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM53_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM53_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM53_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM53_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM53_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM53_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM53_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM53_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM53_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM53_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM53_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM53_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM53_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM53_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM53_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM53_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM53_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM53_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM53_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM53_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM53_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM53_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM53_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM53_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM53_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM53_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM53_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM53_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM53_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM53_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM53_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM53_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM53_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM53_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM53_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM53_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM53_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM53_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM53_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM53_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM53_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM53_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM53_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM53_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM53_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM53_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(53), SSRA=>'0', WEA=>wea , DOA=>DOvecA(53), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(53), SSRb=>'0', WEb=>'0', DOb=>DOvecB(53), DOPb=>open);

RAM54 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM54_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM54_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM54_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM54_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM54_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM54_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM54_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM54_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM54_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM54_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM54_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM54_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM54_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM54_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM54_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM54_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM54_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM54_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM54_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM54_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM54_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM54_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM54_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM54_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM54_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM54_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM54_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM54_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM54_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM54_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM54_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM54_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM54_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM54_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM54_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM54_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM54_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM54_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM54_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM54_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM54_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM54_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM54_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM54_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM54_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM54_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM54_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM54_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM54_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM54_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM54_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM54_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM54_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM54_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM54_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM54_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM54_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM54_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM54_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM54_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM54_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM54_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM54_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM54_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(54), SSRA=>'0', WEA=>wea , DOA=>DOvecA(54), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(54), SSRb=>'0', WEb=>'0', DOb=>DOvecB(54), DOPb=>open);

RAM55 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM55_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM55_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM55_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM55_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM55_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM55_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM55_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM55_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM55_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM55_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM55_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM55_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM55_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM55_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM55_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM55_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM55_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM55_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM55_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM55_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM55_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM55_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM55_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM55_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM55_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM55_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM55_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM55_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM55_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM55_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM55_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM55_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM55_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM55_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM55_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM55_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM55_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM55_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM55_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM55_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM55_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM55_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM55_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM55_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM55_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM55_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM55_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM55_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM55_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM55_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM55_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM55_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM55_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM55_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM55_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM55_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM55_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM55_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM55_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM55_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM55_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM55_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM55_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM55_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(55), SSRA=>'0', WEA=>wea , DOA=>DOvecA(55), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(55), SSRb=>'0', WEb=>'0', DOb=>DOvecB(55), DOPb=>open);

RAM56 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM56_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM56_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM56_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM56_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM56_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM56_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM56_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM56_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM56_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM56_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM56_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM56_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM56_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM56_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM56_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM56_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM56_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM56_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM56_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM56_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM56_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM56_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM56_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM56_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM56_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM56_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM56_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM56_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM56_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM56_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM56_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM56_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM56_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM56_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM56_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM56_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM56_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM56_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM56_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM56_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM56_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM56_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM56_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM56_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM56_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM56_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM56_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM56_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM56_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM56_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM56_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM56_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM56_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM56_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM56_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM56_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM56_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM56_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM56_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM56_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM56_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM56_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM56_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM56_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(56), SSRA=>'0', WEA=>wea , DOA=>DOvecA(56), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(56), SSRb=>'0', WEb=>'0', DOb=>DOvecB(56), DOPb=>open);

RAM57 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM57_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM57_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM57_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM57_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM57_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM57_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM57_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM57_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM57_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM57_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM57_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM57_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM57_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM57_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM57_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM57_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM57_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM57_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM57_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM57_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM57_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM57_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM57_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM57_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM57_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM57_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM57_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM57_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM57_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM57_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM57_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM57_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM57_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM57_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM57_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM57_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM57_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM57_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM57_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM57_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM57_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM57_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM57_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM57_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM57_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM57_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM57_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM57_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM57_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM57_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM57_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM57_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM57_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM57_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM57_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM57_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM57_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM57_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM57_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM57_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM57_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM57_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM57_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM57_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(57), SSRA=>'0', WEA=>wea , DOA=>DOvecA(57), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(57), SSRb=>'0', WEb=>'0', DOb=>DOvecB(57), DOPb=>open);

RAM58 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM58_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM58_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM58_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM58_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM58_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM58_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM58_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM58_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM58_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM58_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM58_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM58_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM58_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM58_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM58_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM58_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM58_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM58_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM58_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM58_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM58_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM58_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM58_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM58_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM58_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM58_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM58_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM58_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM58_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM58_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM58_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM58_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM58_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM58_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM58_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM58_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM58_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM58_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM58_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM58_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM58_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM58_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM58_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM58_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM58_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM58_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM58_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM58_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM58_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM58_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM58_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM58_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM58_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM58_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM58_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM58_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM58_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM58_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM58_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM58_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM58_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM58_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM58_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM58_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(58), SSRA=>'0', WEA=>wea , DOA=>DOvecA(58), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(58), SSRb=>'0', WEb=>'0', DOb=>DOvecB(58), DOPb=>open);

RAM59 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM59_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM59_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM59_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM59_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM59_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM59_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM59_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM59_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM59_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM59_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM59_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM59_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM59_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM59_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM59_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM59_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM59_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM59_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM59_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM59_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM59_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM59_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM59_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM59_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM59_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM59_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM59_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM59_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM59_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM59_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM59_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM59_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM59_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM59_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM59_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM59_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM59_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM59_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM59_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM59_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM59_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM59_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM59_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM59_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM59_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM59_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM59_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM59_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM59_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM59_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM59_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM59_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM59_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM59_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM59_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM59_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM59_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM59_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM59_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM59_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM59_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM59_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM59_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM59_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(59), SSRA=>'0', WEA=>wea , DOA=>DOvecA(59), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(59), SSRb=>'0', WEb=>'0', DOb=>DOvecB(59), DOPb=>open);

RAM60 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM60_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM60_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM60_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM60_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM60_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM60_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM60_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM60_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM60_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM60_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM60_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM60_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM60_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM60_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM60_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM60_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM60_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM60_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM60_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM60_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM60_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM60_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM60_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM60_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM60_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM60_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM60_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM60_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM60_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM60_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM60_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM60_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM60_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM60_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM60_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM60_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM60_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM60_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM60_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM60_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM60_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM60_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM60_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM60_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM60_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM60_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM60_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM60_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM60_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM60_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM60_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM60_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM60_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM60_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM60_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM60_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM60_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM60_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM60_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM60_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM60_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM60_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM60_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM60_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(60), SSRA=>'0', WEA=>wea , DOA=>DOvecA(60), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(60), SSRb=>'0', WEb=>'0', DOb=>DOvecB(60), DOPb=>open);

RAM61 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM61_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM61_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM61_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM61_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM61_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM61_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM61_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM61_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM61_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM61_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM61_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM61_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM61_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM61_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM61_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM61_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM61_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM61_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM61_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM61_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM61_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM61_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM61_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM61_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM61_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM61_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM61_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM61_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM61_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM61_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM61_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM61_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM61_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM61_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM61_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM61_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM61_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM61_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM61_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM61_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM61_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM61_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM61_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM61_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM61_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM61_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM61_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM61_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM61_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM61_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM61_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM61_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM61_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM61_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM61_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM61_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM61_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM61_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM61_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM61_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM61_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM61_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM61_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM61_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(61), SSRA=>'0', WEA=>wea , DOA=>DOvecA(61), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(61), SSRb=>'0', WEb=>'0', DOb=>DOvecB(61), DOPb=>open);

RAM62 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM62_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM62_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM62_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM62_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM62_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM62_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM62_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM62_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM62_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM62_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM62_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM62_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM62_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM62_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM62_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM62_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM62_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM62_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM62_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM62_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM62_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM62_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM62_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM62_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM62_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM62_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM62_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM62_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM62_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM62_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM62_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM62_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM62_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM62_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM62_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM62_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM62_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM62_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM62_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM62_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM62_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM62_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM62_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM62_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM62_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM62_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM62_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM62_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM62_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM62_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM62_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM62_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM62_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM62_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM62_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM62_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM62_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM62_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM62_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM62_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM62_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM62_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM62_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM62_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(62), SSRA=>'0', WEA=>wea , DOA=>DOvecA(62), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(62), SSRb=>'0', WEb=>'0', DOb=>DOvecB(62), DOPb=>open);

RAM63 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM63_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM63_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM63_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM63_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM63_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM63_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM63_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM63_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM63_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM63_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM63_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM63_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM63_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM63_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM63_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM63_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM63_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM63_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM63_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM63_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM63_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM63_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM63_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM63_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM63_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM63_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM63_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM63_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM63_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM63_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM63_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM63_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM63_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM63_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM63_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM63_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM63_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM63_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM63_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM63_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM63_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM63_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM63_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM63_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM63_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM63_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM63_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM63_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM63_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM63_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM63_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM63_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM63_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM63_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM63_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM63_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM63_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM63_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM63_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM63_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM63_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM63_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM63_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM63_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(63), SSRA=>'0', WEA=>wea , DOA=>DOvecA(63), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(63), SSRb=>'0', WEb=>'0', DOb=>DOvecB(63), DOPb=>open);

RAM64 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM64_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM64_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM64_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM64_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM64_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM64_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM64_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM64_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM64_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM64_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM64_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM64_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM64_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM64_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM64_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM64_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM64_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM64_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM64_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM64_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM64_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM64_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM64_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM64_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM64_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM64_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM64_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM64_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM64_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM64_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM64_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM64_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM64_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM64_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM64_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM64_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM64_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM64_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM64_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM64_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM64_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM64_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM64_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM64_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM64_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM64_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM64_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM64_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM64_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM64_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM64_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM64_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM64_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM64_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM64_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM64_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM64_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM64_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM64_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM64_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM64_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM64_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM64_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM64_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(64), SSRA=>'0', WEA=>wea , DOA=>DOvecA(64), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(64), SSRb=>'0', WEb=>'0', DOb=>DOvecB(64), DOPb=>open);

RAM65 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM65_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM65_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM65_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM65_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM65_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM65_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM65_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM65_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM65_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM65_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM65_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM65_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM65_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM65_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM65_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM65_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM65_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM65_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM65_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM65_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM65_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM65_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM65_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM65_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM65_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM65_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM65_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM65_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM65_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM65_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM65_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM65_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM65_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM65_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM65_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM65_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM65_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM65_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM65_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM65_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM65_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM65_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM65_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM65_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM65_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM65_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM65_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM65_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM65_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM65_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM65_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM65_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM65_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM65_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM65_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM65_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM65_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM65_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM65_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM65_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM65_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM65_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM65_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM65_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(65), SSRA=>'0', WEA=>wea , DOA=>DOvecA(65), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(65), SSRb=>'0', WEb=>'0', DOb=>DOvecB(65), DOPb=>open);

RAM66 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM66_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM66_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM66_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM66_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM66_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM66_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM66_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM66_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM66_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM66_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM66_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM66_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM66_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM66_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM66_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM66_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM66_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM66_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM66_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM66_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM66_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM66_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM66_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM66_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM66_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM66_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM66_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM66_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM66_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM66_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM66_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM66_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM66_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM66_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM66_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM66_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM66_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM66_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM66_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM66_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM66_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM66_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM66_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM66_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM66_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM66_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM66_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM66_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM66_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM66_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM66_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM66_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM66_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM66_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM66_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM66_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM66_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM66_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM66_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM66_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM66_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM66_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM66_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM66_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(66), SSRA=>'0', WEA=>wea , DOA=>DOvecA(66), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(66), SSRb=>'0', WEb=>'0', DOb=>DOvecB(66), DOPb=>open);

RAM67 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM67_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM67_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM67_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM67_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM67_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM67_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM67_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM67_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM67_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM67_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM67_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM67_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM67_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM67_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM67_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM67_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM67_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM67_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM67_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM67_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM67_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM67_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM67_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM67_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM67_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM67_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM67_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM67_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM67_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM67_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM67_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM67_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM67_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM67_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM67_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM67_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM67_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM67_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM67_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM67_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM67_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM67_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM67_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM67_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM67_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM67_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM67_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM67_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM67_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM67_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM67_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM67_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM67_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM67_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM67_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM67_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM67_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM67_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM67_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM67_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM67_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM67_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM67_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM67_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(67), SSRA=>'0', WEA=>wea , DOA=>DOvecA(67), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(67), SSRb=>'0', WEb=>'0', DOb=>DOvecB(67), DOPb=>open);

RAM68 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM68_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM68_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM68_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM68_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM68_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM68_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM68_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM68_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM68_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM68_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM68_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM68_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM68_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM68_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM68_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM68_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM68_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM68_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM68_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM68_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM68_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM68_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM68_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM68_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM68_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM68_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM68_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM68_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM68_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM68_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM68_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM68_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM68_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM68_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM68_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM68_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM68_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM68_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM68_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM68_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM68_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM68_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM68_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM68_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM68_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM68_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM68_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM68_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM68_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM68_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM68_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM68_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM68_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM68_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM68_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM68_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM68_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM68_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM68_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM68_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM68_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM68_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM68_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM68_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(68), SSRA=>'0', WEA=>wea , DOA=>DOvecA(68), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(68), SSRb=>'0', WEb=>'0', DOb=>DOvecB(68), DOPb=>open);

RAM69 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM69_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM69_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM69_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM69_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM69_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM69_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM69_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM69_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM69_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM69_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM69_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM69_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM69_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM69_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM69_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM69_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM69_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM69_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM69_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM69_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM69_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM69_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM69_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM69_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM69_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM69_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM69_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM69_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM69_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM69_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM69_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM69_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM69_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM69_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM69_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM69_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM69_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM69_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM69_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM69_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM69_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM69_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM69_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM69_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM69_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM69_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM69_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM69_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM69_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM69_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM69_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM69_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM69_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM69_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM69_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM69_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM69_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM69_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM69_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM69_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM69_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM69_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM69_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM69_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(69), SSRA=>'0', WEA=>wea , DOA=>DOvecA(69), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(69), SSRb=>'0', WEb=>'0', DOb=>DOvecB(69), DOPb=>open);

RAM70 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM70_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM70_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM70_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM70_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM70_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM70_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM70_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM70_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM70_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM70_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM70_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM70_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM70_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM70_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM70_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM70_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM70_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM70_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM70_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM70_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM70_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM70_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM70_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM70_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM70_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM70_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM70_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM70_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM70_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM70_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM70_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM70_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM70_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM70_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM70_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM70_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM70_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM70_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM70_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM70_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM70_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM70_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM70_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM70_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM70_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM70_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM70_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM70_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM70_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM70_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM70_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM70_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM70_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM70_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM70_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM70_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM70_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM70_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM70_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM70_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM70_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM70_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM70_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM70_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(70), SSRA=>'0', WEA=>wea , DOA=>DOvecA(70), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(70), SSRb=>'0', WEb=>'0', DOb=>DOvecB(70), DOPb=>open);

RAM71 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM71_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM71_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM71_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM71_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM71_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM71_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM71_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM71_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM71_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM71_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM71_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM71_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM71_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM71_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM71_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM71_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM71_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM71_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM71_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM71_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM71_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM71_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM71_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM71_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM71_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM71_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM71_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM71_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM71_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM71_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM71_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM71_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM71_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM71_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM71_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM71_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM71_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM71_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM71_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM71_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM71_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM71_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM71_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM71_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM71_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM71_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM71_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM71_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM71_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM71_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM71_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM71_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM71_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM71_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM71_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM71_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM71_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM71_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM71_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM71_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM71_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM71_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM71_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM71_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(71), SSRA=>'0', WEA=>wea , DOA=>DOvecA(71), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(71), SSRb=>'0', WEb=>'0', DOb=>DOvecB(71), DOPb=>open);

RAM72 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM72_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM72_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM72_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM72_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM72_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM72_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM72_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM72_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM72_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM72_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM72_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM72_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM72_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM72_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM72_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM72_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM72_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM72_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM72_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM72_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM72_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM72_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM72_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM72_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM72_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM72_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM72_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM72_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM72_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM72_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM72_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM72_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM72_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM72_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM72_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM72_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM72_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM72_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM72_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM72_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM72_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM72_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM72_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM72_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM72_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM72_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM72_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM72_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM72_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM72_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM72_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM72_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM72_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM72_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM72_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM72_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM72_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM72_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM72_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM72_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM72_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM72_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM72_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM72_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(72), SSRA=>'0', WEA=>wea , DOA=>DOvecA(72), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(72), SSRb=>'0', WEb=>'0', DOb=>DOvecB(72), DOPb=>open);

RAM73 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM73_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM73_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM73_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM73_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM73_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM73_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM73_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM73_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM73_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM73_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM73_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM73_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM73_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM73_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM73_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM73_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM73_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM73_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM73_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM73_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM73_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM73_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM73_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM73_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM73_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM73_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM73_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM73_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM73_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM73_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM73_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM73_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM73_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM73_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM73_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM73_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM73_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM73_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM73_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM73_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM73_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM73_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM73_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM73_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM73_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM73_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM73_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM73_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM73_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM73_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM73_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM73_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM73_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM73_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM73_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM73_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM73_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM73_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM73_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM73_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM73_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM73_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM73_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM73_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(73), SSRA=>'0', WEA=>wea , DOA=>DOvecA(73), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(73), SSRb=>'0', WEb=>'0', DOb=>DOvecB(73), DOPb=>open);

RAM74 : RAMB16_S18_S18
generic map (
INIT_00=>C_VGA_C_RAM_VIDEO_RAM74_INIT_00, INIT_01=>C_VGA_C_RAM_VIDEO_RAM74_INIT_01, INIT_02=>C_VGA_C_RAM_VIDEO_RAM74_INIT_02, INIT_03=>C_VGA_C_RAM_VIDEO_RAM74_INIT_03,
INIT_04=>C_VGA_C_RAM_VIDEO_RAM74_INIT_04, INIT_05=>C_VGA_C_RAM_VIDEO_RAM74_INIT_05, INIT_06=>C_VGA_C_RAM_VIDEO_RAM74_INIT_06, INIT_07=>C_VGA_C_RAM_VIDEO_RAM74_INIT_07,
INIT_08=>C_VGA_C_RAM_VIDEO_RAM74_INIT_08, INIT_09=>C_VGA_C_RAM_VIDEO_RAM74_INIT_09, INIT_0a=>C_VGA_C_RAM_VIDEO_RAM74_INIT_0A, INIT_0b=>C_VGA_C_RAM_VIDEO_RAM74_INIT_0B,
INIT_0c=>C_VGA_C_RAM_VIDEO_RAM74_INIT_0C, INIT_0d=>C_VGA_C_RAM_VIDEO_RAM74_INIT_0D, INIT_0e=>C_VGA_C_RAM_VIDEO_RAM74_INIT_0E, INIT_0f=>C_VGA_C_RAM_VIDEO_RAM74_INIT_0F,
INIT_10=>C_VGA_C_RAM_VIDEO_RAM74_INIT_10, INIT_11=>C_VGA_C_RAM_VIDEO_RAM74_INIT_11, INIT_12=>C_VGA_C_RAM_VIDEO_RAM74_INIT_12, INIT_13=>C_VGA_C_RAM_VIDEO_RAM74_INIT_13,
INIT_14=>C_VGA_C_RAM_VIDEO_RAM74_INIT_14, INIT_15=>C_VGA_C_RAM_VIDEO_RAM74_INIT_15, INIT_16=>C_VGA_C_RAM_VIDEO_RAM74_INIT_16, INIT_17=>C_VGA_C_RAM_VIDEO_RAM74_INIT_17,
INIT_18=>C_VGA_C_RAM_VIDEO_RAM74_INIT_18, INIT_19=>C_VGA_C_RAM_VIDEO_RAM74_INIT_19, INIT_1a=>C_VGA_C_RAM_VIDEO_RAM74_INIT_1A, INIT_1b=>C_VGA_C_RAM_VIDEO_RAM74_INIT_1B,
INIT_1c=>C_VGA_C_RAM_VIDEO_RAM74_INIT_1C, INIT_1d=>C_VGA_C_RAM_VIDEO_RAM74_INIT_1D, INIT_1e=>C_VGA_C_RAM_VIDEO_RAM74_INIT_1E, INIT_1f=>C_VGA_C_RAM_VIDEO_RAM74_INIT_1F,
INIT_20=>C_VGA_C_RAM_VIDEO_RAM74_INIT_20, INIT_21=>C_VGA_C_RAM_VIDEO_RAM74_INIT_21, INIT_22=>C_VGA_C_RAM_VIDEO_RAM74_INIT_22, INIT_23=>C_VGA_C_RAM_VIDEO_RAM74_INIT_23,
INIT_24=>C_VGA_C_RAM_VIDEO_RAM74_INIT_24, INIT_25=>C_VGA_C_RAM_VIDEO_RAM74_INIT_25, INIT_26=>C_VGA_C_RAM_VIDEO_RAM74_INIT_26, INIT_27=>C_VGA_C_RAM_VIDEO_RAM74_INIT_27,
INIT_28=>C_VGA_C_RAM_VIDEO_RAM74_INIT_28, INIT_29=>C_VGA_C_RAM_VIDEO_RAM74_INIT_29, INIT_2a=>C_VGA_C_RAM_VIDEO_RAM74_INIT_2A, INIT_2b=>C_VGA_C_RAM_VIDEO_RAM74_INIT_2B,
INIT_2c=>C_VGA_C_RAM_VIDEO_RAM74_INIT_2C, INIT_2d=>C_VGA_C_RAM_VIDEO_RAM74_INIT_2D, INIT_2e=>C_VGA_C_RAM_VIDEO_RAM74_INIT_2E, INIT_2f=>C_VGA_C_RAM_VIDEO_RAM74_INIT_2F,
INIT_30=>C_VGA_C_RAM_VIDEO_RAM74_INIT_30, INIT_31=>C_VGA_C_RAM_VIDEO_RAM74_INIT_31, INIT_32=>C_VGA_C_RAM_VIDEO_RAM74_INIT_32, INIT_33=>C_VGA_C_RAM_VIDEO_RAM74_INIT_33,
INIT_34=>C_VGA_C_RAM_VIDEO_RAM74_INIT_34, INIT_35=>C_VGA_C_RAM_VIDEO_RAM74_INIT_35, INIT_36=>C_VGA_C_RAM_VIDEO_RAM74_INIT_36, INIT_37=>C_VGA_C_RAM_VIDEO_RAM74_INIT_37,
INIT_38=>C_VGA_C_RAM_VIDEO_RAM74_INIT_38, INIT_39=>C_VGA_C_RAM_VIDEO_RAM74_INIT_39, INIT_3a=>C_VGA_C_RAM_VIDEO_RAM74_INIT_3A, INIT_3b=>C_VGA_C_RAM_VIDEO_RAM74_INIT_3B,
INIT_3c=>C_VGA_C_RAM_VIDEO_RAM74_INIT_3C, INIT_3d=>C_VGA_C_RAM_VIDEO_RAM74_INIT_3D, INIT_3e=>C_VGA_C_RAM_VIDEO_RAM74_INIT_3E, INIT_3f=>C_VGA_C_RAM_VIDEO_RAM74_INIT_3F)
port map (ADDRA=>std_logic_vector(addra(9 downto 0)), CLKA=> CLKA, DIA=> std_logic_vector(dia), DIPA=>"00", ENA=>ena(74), SSRA=>'0', WEA=>wea , DOA=>DOvecA(74), DOPA=>open,
ADDRb=>std_logic_vector(addrb(9 downto 0)), CLKb=> CLKb, DIb=> X"0000", DIPb=>"00", ENb=>enb(74), SSRb=>'0', WEb=>'0', DOb=>DOvecB(74), DOPb=>open);

end BEHAVIORAL;
