library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
Library UNISIM;
use UNISIM.vcomponents.all;
    
RAMB36E1_inst : RAMB36E1
generic map (
-- Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE"
                RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
-- Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
                SIM_COLLISION_CHECK => "ALL",
-- DOA_REG, DOB_REG: Optional output register (0 or 1)
                DOA_REG => 0,
                DOB_REG => 0,
                EN_ECC_READ => FALSE,
                EN_ECC_WRITE => FALSE,
-- INITP_00 to INITP_0F: Initial contents of the parity memory array
                INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_0a => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_0b => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_0c => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_0d => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_0e => X"0000000000000000000000000000000000000000000000000000000000000000",
                INITP_0f => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_00 to INIT_7F: Initial contents of the data memory array
                INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_0a => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_0b => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_0c => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_0d => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_0e => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_0f => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1a => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1b => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1c => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1d => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1e => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1f => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2a => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2b => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2c => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2d => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2e => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2f => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3a => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3b => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3c => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3d => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3e => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3f => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_4a => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_4b => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_4c => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_4d => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_4e => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_4f => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_5a => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_5b => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_5c => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_5d => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_5e => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_5f => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_6a => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_6b => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_6c => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_6d => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_6e => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_6f => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_7a => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_7b => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_7c => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_7d => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_7e => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_7f => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_A, INIT_B: Initial values on output ports
                INIT_A => X"000000000",
                INIT_B => X"000000000",
-- Initialization File: RAM initialization
                file INIT_FILE => "NONE",
-- RAM Mode: "SDP" or "TDP"
                RAM_MODE => "TDP",
-- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
                RAM_EXTENSION_A => "NONE",
                RAM_EXTENSION_B => "NONE",
-- READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
                READ_WIDTH_A => 8, -- 0-72
                READ_WIDTH_B => 0, -- 0-36
                WRITE_WIDTH_A => 0, -- 0-36
                WRITE_WIDTH_B => 0, -- 0-72
-- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
                RSTREG_PRIORITY_A => "RSTREG",
                RSTREG_PRIORITY_B => "RSTREG",
-- SRVAL_A, SRVAL_B: Set/reset value for output
                SRVAL_A => X"000000000",
                SRVAL_B => X"000000000",
-- Simulation Device: Must be set to "7SERIES" for simulation behavior
                SIM_DEVICE => "7SERIES",
-- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
                WRITE_MODE_A => "WRITE_FIRST",
                WRITE_MODE_B => "WRITE_FIRST"
            )
port
map
(
)

entity RAM_VIDEO is
  port ( 
    clk  : in    std_logic;   
    addr : in    unsigned (16 downto 0); 
    do   : out   unsigned(23 downto 0)
    );
end RAM_VIDEO;

architecture Behavioral of RAM_VIDEO is
  subtype mot is unsigned( 23 downto 0 );
  type zone_memoire is array (natural range 0 to 640*480/4-1) of mot;
  signal ROM: zone_memoire :=(
--   0 => x"ffffff",
--   1 => x"ffff0f",
--   2 => x"ffffff",
--   3 => x"ffffff",
--   4 => x"ffffff",
--   5 => x"ffffff",
--   6 => x"ffffff",
--   7 => x"ffffff",
--   8 => x"fffff0",
   others => x"000000"
    );
begin
  process(CLK)
  begin 
    if (CLK'event AND CLK='1') then
      do <= ROM(to_integer(addr));
    end if;
  end process;
end Behavioral;
